magic
tech scmos
timestamp 1699617317
<< nwell >>
rect -21 11 20 29
<< polysilicon >>
rect -3 23 0 26
rect -3 3 0 18
rect -3 -16 0 -1
rect -3 -25 0 -21
<< ndiffusion >>
rect -6 -21 -3 -16
rect 0 -21 4 -16
<< pdiffusion >>
rect -7 18 -3 23
rect 0 18 4 23
rect 8 18 10 23
<< metal1 >>
rect -21 29 -8 33
rect -4 29 20 33
rect -11 23 -8 29
rect -6 -1 -4 3
rect 5 -16 8 18
rect -11 -28 -7 -21
rect -21 -34 21 -28
<< ntransistor >>
rect -3 -21 0 -16
<< ptransistor >>
rect -3 18 0 23
<< polycontact >>
rect -4 -1 0 3
<< ndcontact >>
rect -11 -21 -6 -16
rect 4 -21 8 -16
<< pdcontact >>
rect -11 18 -7 23
rect 4 18 8 23
<< nsubstratencontact >>
rect -8 29 -4 33
<< labels >>
rlabel metal1 -5 1 -5 1 1 A
rlabel metal1 6 0 6 0 1 out
rlabel metal1 2 31 2 31 5 vdd
rlabel metal1 -3 -31 -3 -31 1 gnd
<< end >>
