* SPICE3 file created from adder_subtractor.ext - technology: scmos

.include TSMC_180nm.txt


.param SUPPLY = 1
.param LAMBDA = 0.18u

.param width_P=8*LAMBDA
.param  width_N = 4*LAMBDA
.global gnd vdd
.option scale=0.09u

Vdd vdd gnd 'SUPPLY'


* Va3 A1 gnd PULSE(1.8 0 400ns 100ps 100ps 400ns 800ns)
* * Va2 a2 gnd PULSE(0 1.8 400ns 100ps 100ps 400ns 800ns)
* * Va1 A1 gnd PULSE(1.8 0 400ns 100ps 100ps 400ns 800ns)
* Va0 A0 gnd PULSE(0 1.8 100ns 100ps 100ps 200ns 400ns)


* Vb0 B1 gnd PULSE(0 1.8 100ns 100ps 100ps 200ns 400ns)
* * Va2 a2 gnd PULSE(0 1.8 400ns 100ps 100ps 400ns 800ns)
* * Va1 A1 gnd PULSE(1.8 0 400ns 100ps 100ps 400ns 800ns)
* Vb3 B0 gnd PULSE(1.8 0 400ns 100ps 100ps 400ns 800ns)


VE M 0 DC 1V

Va3 a3 0 DC 1V
Va2 a2 0 DC 1V
Va1 a1 0 DC 1V
Va0 a0 0 DC 1V
* even if the inputs are 1 , it will consider 1.8 because of supply ( MOSFETS ) ON AND OFF 

Vb3 b3 0 DC 1V
Vb2 b2 0 DC 1V
Vb1 b1 0 DC 0V
Vb0 b0 0 DC 1V


.option scale=1u


M1000 a_n1544_n689# C2 vdd w_n1536_n653# CMOSP w=5 l=2
+  ad=30 pd=22 as=2880 ps=1808
M1001 a_n579_n673# a_n894_n765# a_n579_n706# Gnd CMOSN w=9 l=3
+  ad=72 pd=34 as=72 ps=34
M1002 a_n1732_n679# a_n1749_n693# a_n1720_n679# w_n1741_n657# CMOSP w=5 l=2
+  ad=85 pd=64 as=55 ps=42
M1003 a_n2258_n792# a_n2316_n755# gnd Gnd CMOSN w=5 l=3
+  ad=40 pd=26 as=2000 ps=1288
M1004 a_n155_n657# a_n44_n522# B0 Gnd CMOSN w=5 l=2
+  ad=58 pd=44 as=23 ps=20
M1005 a_n152_n734# A0 vdd w_n167_n737# CMOSP w=7 l=3
+  ad=56 pd=30 as=0 ps=0
M1006 a_64_n670# a_n153_n674# vdd w_43_n648# CMOSP w=5 l=2
+  ad=55 pd=42 as=0 ps=0
M1007 a_n155_n657# M a_n15_n508# Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=50 ps=42
M1008 a_n1731_n772# A2 gnd Gnd CMOSN w=9 l=3
+  ad=72 pd=34 as=0 ps=0
M1009 a_n955_n651# M a_n815_n502# Gnd CMOSN w=5 l=2
+  ad=58 pd=44 as=50 ps=42
M1010 a_3_n767# a_n153_n674# gnd Gnd CMOSN w=9 l=3
+  ad=72 pd=34 as=0 ps=0
M1011 a_n152_n734# a_n155_n657# a_n152_n767# Gnd CMOSN w=9 l=3
+  ad=72 pd=34 as=72 ps=34
M1012 a_n1305_n787# a_n1518_n776# vdd w_n1295_n688# CMOSP w=7 l=3
+  ad=56 pd=30 as=0 ps=0
M1013 vdd C2 a_n1576_n739# w_n1591_n742# CMOSP w=7 l=3
+  ad=0 pd=0 as=56 ps=30
M1014 C2 a_n579_n673# a_n522_n801# Gnd CMOSN w=9 l=3
+  ad=72 pd=34 as=72 ps=34
M1015 a_n153_n674# a_n155_n657# A0 w_n162_n652# CMOSP w=5 l=2
+  ad=85 pd=64 as=25 ps=20
M1016 a_n44_n522# M gnd Gnd CMOSN w=5 l=2
+  ad=28 pd=22 as=0 ps=0
M1017 a_n2041_n828# a_n2045_n803# gnd Gnd CMOSN w=9 l=3
+  ad=72 pd=34 as=0 ps=0
M1018 a_n2489_n709# a_n2474_n678# vdd w_n2481_n673# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1019 S2 a_n1544_n689# a_n1732_n679# Gnd CMOSN w=5 l=2
+  ad=58 pd=44 as=81 ps=64
M1020 vdd a_n2098_n700# carry w_n2056_n798# CMOSP w=7 l=3
+  ad=0 pd=0 as=56 ps=30
M1021 a_n1544_n689# C2 gnd Gnd CMOSN w=5 l=2
+  ad=28 pd=22 as=0 ps=0
M1022 a_n797_n728# a_n953_n668# vdd w_n812_n731# CMOSP w=7 l=3
+  ad=56 pd=30 as=0 ps=0
M1023 a_n1594_n513# B2 gnd Gnd CMOSN w=5 l=2
+  ad=50 pd=42 as=0 ps=0
M1024 a_n1732_n679# a_n1734_n662# a_n1720_n679# Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=50 ps=42
M1025 a_n2098_n733# a_n2413_n792# gnd Gnd CMOSN w=9 l=3
+  ad=72 pd=34 as=0 ps=0
M1026 a_64_n670# a_n153_n674# gnd Gnd CMOSN w=5 l=2
+  ad=50 pd=42 as=0 ps=0
M1027 a_n1734_n662# M a_n1594_n513# Gnd CMOSN w=5 l=2
+  ad=58 pd=44 as=0 ps=0
M1028 a_n15_n508# B0 vdd w_n36_n486# CMOSP w=5 l=2
+  ad=55 pd=42 as=0 ps=0
M1029 S3 C3 a_n2472_n695# w_n2276_n669# CMOSP w=5 l=2
+  ad=60 pd=44 as=85 ps=64
M1030 a_n1518_n776# a_n1576_n739# gnd Gnd CMOSN w=5 l=3
+  ad=40 pd=26 as=0 ps=0
M1031 a_n1305_n787# a_n1518_n776# a_n1280_n718# Gnd CMOSN w=9 l=3
+  ad=72 pd=34 as=72 ps=34
M1032 a_n1734_n662# M B2 w_n1615_n491# CMOSP w=5 l=2
+  ad=60 pd=44 as=25 ps=20
M1033 a_n2255_n691# a_n2472_n695# gnd Gnd CMOSN w=5 l=2
+  ad=50 pd=42 as=0 ps=0
M1034 vdd a_61_n771# a_274_n782# w_284_n683# CMOSP w=7 l=3
+  ad=0 pd=0 as=56 ps=30
M1035 a_n2460_n695# A3 vdd w_n2481_n673# CMOSP w=5 l=2
+  ad=55 pd=42 as=0 ps=0
M1036 C3 a_n1358_n684# a_n1301_n812# Gnd CMOSN w=9 l=3
+  ad=72 pd=34 as=72 ps=34
M1037 a_n1623_n527# M vdd w_n1615_n491# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1038 S3 C3 a_n2255_n691# Gnd CMOSN w=5 l=2
+  ad=58 pd=44 as=0 ps=0
M1039 vdd a_n1673_n776# a_n1358_n684# w_n1373_n687# CMOSP w=7 l=3
+  ad=0 pd=0 as=56 ps=30
M1040 a_n153_n674# a_n170_n688# A0 Gnd CMOSN w=5 l=2
+  ad=81 pd=64 as=23 ps=20
M1041 a_n952_n728# a_n955_n651# a_n952_n761# Gnd CMOSN w=9 l=3
+  ad=72 pd=34 as=72 ps=34
M1042 a_n2413_n792# a_n2471_n755# vdd vdd CMOSP w=5 l=3
+  ad=50 pd=30 as=0 ps=0
M1043 a_n2489_n709# a_n2474_n678# gnd Gnd CMOSN w=5 l=2
+  ad=28 pd=22 as=0 ps=0
M1044 a_n2471_n788# A3 gnd Gnd CMOSN w=9 l=3
+  ad=72 pd=34 as=0 ps=0
M1045 S2 a_n1544_n689# a_n1515_n675# w_n1536_n653# CMOSP w=5 l=2
+  ad=60 pd=44 as=55 ps=42
M1046 vdd a_n739_n765# a_n526_n776# w_n516_n677# CMOSP w=7 l=3
+  ad=0 pd=0 as=56 ps=30
M1047 S0 M a_n153_n674# w_43_n648# CMOSP w=5 l=2
+  ad=60 pd=44 as=0 ps=0
M1048 a_n2316_n788# a_n2472_n695# gnd Gnd CMOSN w=9 l=3
+  ad=72 pd=34 as=0 ps=0
M1049 a_n2460_n695# A3 gnd Gnd CMOSN w=5 l=2
+  ad=50 pd=42 as=0 ps=0
M1050 vdd a_n2474_n678# a_n2471_n755# w_n2486_n758# CMOSP w=7 l=3
+  ad=0 pd=0 as=56 ps=30
M1051 a_n141_n674# A0 vdd w_n162_n652# CMOSP w=5 l=2
+  ad=55 pd=42 as=0 ps=0
M1052 C2 a_n526_n776# vdd w_n537_n771# CMOSP w=7 l=3
+  ad=56 pd=30 as=0 ps=0
M1053 a_n153_n674# a_n170_n688# a_n141_n674# w_n162_n652# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1054 S0 a_35_n684# a_64_n670# w_43_n648# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1055 a_n15_n508# B0 gnd Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1056 a_n2474_n678# M B3 w_n2355_n507# CMOSP w=5 l=2
+  ad=60 pd=44 as=25 ps=20
M1057 S2 C2 a_n1515_n675# Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=50 ps=42
M1058 a_n1734_n662# a_n1623_n527# B2 Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=23 ps=20
M1059 a_221_n712# a_n94_n771# gnd Gnd CMOSN w=9 l=3
+  ad=72 pd=34 as=0 ps=0
M1060 a_n2363_n543# M vdd w_n2355_n507# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1061 vdd a_n2413_n792# a_n2098_n700# w_n2113_n703# CMOSP w=7 l=3
+  ad=0 pd=0 as=56 ps=30
M1062 vdd C3 a_n2316_n755# w_n2331_n758# CMOSP w=7 l=3
+  ad=0 pd=0 as=56 ps=30
M1063 S0 a_35_n684# a_n153_n674# Gnd CMOSN w=5 l=2
+  ad=58 pd=44 as=0 ps=0
M1064 a_n1623_n527# M gnd Gnd CMOSN w=5 l=2
+  ad=28 pd=22 as=0 ps=0
M1065 a_n2255_n691# a_n2472_n695# vdd w_n2276_n669# CMOSP w=5 l=2
+  ad=55 pd=42 as=0 ps=0
M1066 a_n1576_n739# C2 a_n1576_n772# Gnd CMOSN w=9 l=3
+  ad=72 pd=34 as=72 ps=34
M1067 S3 a_n2284_n705# a_n2255_n691# w_n2276_n669# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1068 a_61_n771# a_3_n734# gnd Gnd CMOSN w=5 l=3
+  ad=40 pd=26 as=0 ps=0
M1069 a_n739_n765# a_n797_n728# vdd vdd CMOSP w=5 l=3
+  ad=50 pd=30 as=0 ps=0
M1070 a_n141_n674# A0 gnd Gnd CMOSN w=5 l=2
+  ad=50 pd=42 as=0 ps=0
M1071 a_n2284_n705# C3 gnd Gnd CMOSN w=5 l=2
+  ad=28 pd=22 as=0 ps=0
M1072 a_n797_n761# a_n953_n668# gnd Gnd CMOSN w=9 l=3
+  ad=72 pd=34 as=0 ps=0
M1073 a_n1673_n776# a_n1731_n739# gnd Gnd CMOSN w=5 l=3
+  ad=40 pd=26 as=0 ps=0
M1074 a_n2045_n803# a_n2258_n792# vdd w_n2035_n704# CMOSP w=7 l=3
+  ad=56 pd=30 as=0 ps=0
M1075 a_274_n782# a_61_n771# vdd w_284_n683# CMOSP w=7 l=3
+  ad=0 pd=0 as=0 ps=0
M1076 a_n153_n674# a_n155_n657# a_n141_n674# Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1077 vdd a_n1734_n662# a_n1731_n739# w_n1746_n742# CMOSP w=7 l=3
+  ad=0 pd=0 as=56 ps=30
M1078 S0 M a_64_n670# Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1079 a_n2045_n803# a_n2258_n792# a_n2020_n734# Gnd CMOSN w=9 l=3
+  ad=72 pd=34 as=72 ps=34
M1080 a_n1358_n684# a_n1673_n776# vdd w_n1373_n687# CMOSP w=7 l=3
+  ad=0 pd=0 as=0 ps=0
M1081 vdd M a_3_n734# w_n12_n737# CMOSP w=7 l=3
+  ad=0 pd=0 as=56 ps=30
M1082 a_n170_n688# a_n155_n657# vdd w_n162_n652# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1083 a_n952_n728# A1 vdd w_n967_n731# CMOSP w=7 l=3
+  ad=56 pd=30 as=0 ps=0
M1084 vdd a_221_n679# C1 w_263_n777# CMOSP w=7 l=3
+  ad=0 pd=0 as=56 ps=30
M1085 a_n2474_n678# a_n2363_n543# B3 Gnd CMOSN w=5 l=2
+  ad=58 pd=44 as=23 ps=20
M1086 a_n2363_n543# M gnd Gnd CMOSN w=5 l=2
+  ad=28 pd=22 as=0 ps=0
M1087 a_n953_n668# a_n955_n651# A1 w_n962_n646# CMOSP w=5 l=2
+  ad=85 pd=64 as=25 ps=20
M1088 a_274_n782# a_61_n771# a_299_n713# Gnd CMOSN w=9 l=3
+  ad=72 pd=34 as=72 ps=34
M1089 a_n2334_n529# B3 vdd w_n2355_n507# CMOSP w=5 l=2
+  ad=55 pd=42 as=0 ps=0
M1090 a_n970_n682# a_n955_n651# vdd w_n962_n646# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1091 a_n94_n771# a_n152_n734# vdd vdd CMOSP w=5 l=3
+  ad=50 pd=30 as=0 ps=0
M1092 a_n2474_n678# a_n2363_n543# a_n2334_n529# w_n2355_n507# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1093 a_278_n807# a_274_n782# gnd Gnd CMOSN w=9 l=3
+  ad=72 pd=34 as=0 ps=0
M1094 vdd a_n94_n771# a_221_n679# w_206_n682# CMOSP w=7 l=3
+  ad=0 pd=0 as=56 ps=30
M1095 a_n170_n688# a_n155_n657# gnd Gnd CMOSN w=5 l=2
+  ad=28 pd=22 as=0 ps=0
M1096 a_n579_n706# a_n894_n765# gnd Gnd CMOSN w=9 l=3
+  ad=0 pd=0 as=0 ps=0
M1097 a_n2284_n705# C3 vdd w_n2276_n669# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1098 vdd a_n894_n765# a_n579_n673# w_n594_n676# CMOSP w=7 l=3
+  ad=0 pd=0 as=56 ps=30
M1099 a_n953_n668# a_n970_n682# A1 Gnd CMOSN w=5 l=2
+  ad=81 pd=64 as=23 ps=20
M1100 a_n152_n767# A0 gnd Gnd CMOSN w=9 l=3
+  ad=0 pd=0 as=0 ps=0
M1101 a_n501_n707# a_n739_n765# gnd Gnd CMOSN w=9 l=3
+  ad=72 pd=34 as=0 ps=0
M1102 S1 a_n765_n678# a_n736_n664# w_n757_n642# CMOSP w=5 l=2
+  ad=60 pd=44 as=55 ps=42
M1103 a_n970_n682# a_n955_n651# gnd Gnd CMOSN w=5 l=2
+  ad=28 pd=22 as=0 ps=0
M1104 a_n1576_n739# a_n1732_n679# vdd w_n1591_n742# CMOSP w=7 l=3
+  ad=0 pd=0 as=0 ps=0
M1105 a_n894_n765# a_n952_n728# vdd vdd CMOSP w=5 l=3
+  ad=50 pd=30 as=0 ps=0
M1106 a_n522_n801# a_n526_n776# gnd Gnd CMOSN w=9 l=3
+  ad=0 pd=0 as=0 ps=0
M1107 a_n815_n502# B1 vdd w_n836_n480# CMOSP w=5 l=2
+  ad=55 pd=42 as=0 ps=0
M1108 carry a_n2045_n803# vdd w_n2056_n798# CMOSP w=7 l=3
+  ad=0 pd=0 as=0 ps=0
M1109 a_n2413_n792# a_n2471_n755# gnd Gnd CMOSN w=5 l=3
+  ad=40 pd=26 as=0 ps=0
M1110 a_n2098_n700# a_n2413_n792# a_n2098_n733# Gnd CMOSN w=9 l=3
+  ad=72 pd=34 as=0 ps=0
M1111 a_n2334_n529# B3 gnd Gnd CMOSN w=5 l=2
+  ad=50 pd=42 as=0 ps=0
M1112 S1 C1 a_n953_n668# w_n757_n642# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1113 a_3_n734# a_n153_n674# vdd w_n12_n737# CMOSP w=7 l=3
+  ad=0 pd=0 as=0 ps=0
M1114 vdd a_n155_n657# a_n152_n734# w_n167_n737# CMOSP w=7 l=3
+  ad=0 pd=0 as=0 ps=0
M1115 a_n941_n668# A1 vdd w_n962_n646# CMOSP w=5 l=2
+  ad=55 pd=42 as=0 ps=0
M1116 a_n1731_n739# a_n1734_n662# a_n1731_n772# Gnd CMOSN w=9 l=3
+  ad=72 pd=34 as=0 ps=0
M1117 a_n1280_n718# a_n1518_n776# gnd Gnd CMOSN w=9 l=3
+  ad=0 pd=0 as=0 ps=0
M1118 a_n2474_n678# M a_n2334_n529# Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1119 a_n765_n678# C1 vdd w_n757_n642# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1120 S1 C1 a_n736_n664# Gnd CMOSN w=5 l=2
+  ad=58 pd=44 as=50 ps=42
M1121 vdd a_n1518_n776# a_n1305_n787# w_n1295_n688# CMOSP w=7 l=3
+  ad=0 pd=0 as=0 ps=0
M1122 a_n953_n668# a_n970_n682# a_n941_n668# w_n962_n646# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1123 carry a_n2098_n700# a_n2041_n828# Gnd CMOSN w=9 l=3
+  ad=72 pd=34 as=0 ps=0
M1124 a_n952_n761# A1 gnd Gnd CMOSN w=9 l=3
+  ad=0 pd=0 as=0 ps=0
M1125 a_299_n713# a_61_n771# gnd Gnd CMOSN w=9 l=3
+  ad=0 pd=0 as=0 ps=0
M1126 a_n2258_n792# a_n2316_n755# vdd vdd CMOSP w=5 l=3
+  ad=50 pd=30 as=0 ps=0
M1127 vdd C1 a_n797_n728# w_n812_n731# CMOSP w=7 l=3
+  ad=0 pd=0 as=0 ps=0
M1128 S1 a_n765_n678# a_n953_n668# Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1129 C3 a_n1305_n787# vdd w_n1316_n782# CMOSP w=7 l=3
+  ad=56 pd=30 as=0 ps=0
M1130 a_n941_n668# A1 gnd Gnd CMOSN w=5 l=2
+  ad=50 pd=42 as=0 ps=0
M1131 a_n765_n678# C1 gnd Gnd CMOSN w=5 l=2
+  ad=28 pd=22 as=0 ps=0
M1132 a_n1358_n684# a_n1673_n776# a_n1358_n717# Gnd CMOSN w=9 l=3
+  ad=72 pd=34 as=72 ps=34
M1133 a_n815_n502# B1 gnd Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1134 a_n953_n668# a_n955_n651# a_n941_n668# Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1135 a_n2471_n755# A3 vdd w_n2486_n758# CMOSP w=7 l=3
+  ad=0 pd=0 as=0 ps=0
M1136 a_n2471_n755# a_n2474_n678# a_n2471_n788# Gnd CMOSN w=9 l=3
+  ad=72 pd=34 as=0 ps=0
M1137 a_n526_n776# a_n739_n765# a_n501_n707# Gnd CMOSN w=9 l=3
+  ad=72 pd=34 as=0 ps=0
M1138 a_n955_n651# M B1 w_n836_n480# CMOSP w=5 l=2
+  ad=60 pd=44 as=25 ps=20
M1139 a_n739_n765# a_n797_n728# gnd Gnd CMOSN w=5 l=3
+  ad=40 pd=26 as=0 ps=0
M1140 a_n2472_n695# a_n2474_n678# A3 w_n2481_n673# CMOSP w=5 l=2
+  ad=0 pd=0 as=25 ps=20
M1141 a_n844_n516# M vdd w_n836_n480# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1142 a_221_n679# a_n94_n771# a_221_n712# Gnd CMOSN w=9 l=3
+  ad=72 pd=34 as=0 ps=0
M1143 a_n736_n664# a_n953_n668# vdd w_n757_n642# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1144 a_n1518_n776# a_n1576_n739# vdd vdd CMOSP w=5 l=3
+  ad=50 pd=30 as=0 ps=0
M1145 a_n2316_n755# a_n2472_n695# vdd w_n2331_n758# CMOSP w=7 l=3
+  ad=0 pd=0 as=0 ps=0
M1146 a_n1576_n772# a_n1732_n679# gnd Gnd CMOSN w=9 l=3
+  ad=0 pd=0 as=0 ps=0
M1147 a_n2316_n755# C3 a_n2316_n788# Gnd CMOSN w=9 l=3
+  ad=72 pd=34 as=0 ps=0
M1148 vdd a_n579_n673# C2 w_n537_n771# CMOSP w=7 l=3
+  ad=0 pd=0 as=0 ps=0
M1149 a_n1731_n739# A2 vdd w_n1746_n742# CMOSP w=7 l=3
+  ad=0 pd=0 as=0 ps=0
M1150 a_35_n684# M vdd w_43_n648# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1151 a_n2472_n695# a_n2489_n709# A3 Gnd CMOSN w=5 l=2
+  ad=81 pd=64 as=23 ps=20
M1152 a_n2020_n734# a_n2258_n792# gnd Gnd CMOSN w=9 l=3
+  ad=0 pd=0 as=0 ps=0
M1153 a_n1515_n675# a_n1732_n679# vdd w_n1536_n653# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1154 a_n2098_n700# a_n2413_n792# vdd w_n2113_n703# CMOSP w=7 l=3
+  ad=0 pd=0 as=0 ps=0
M1155 a_n1732_n679# a_n1734_n662# A2 w_n1741_n657# CMOSP w=5 l=2
+  ad=0 pd=0 as=25 ps=20
M1156 a_n736_n664# a_n953_n668# gnd Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1157 a_3_n734# M a_3_n767# Gnd CMOSN w=9 l=3
+  ad=72 pd=34 as=0 ps=0
M1158 a_n94_n771# a_n152_n734# gnd Gnd CMOSN w=5 l=3
+  ad=40 pd=26 as=0 ps=0
M1159 a_n955_n651# a_n844_n516# B1 Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=23 ps=20
M1160 a_n1749_n693# a_n1734_n662# vdd w_n1741_n657# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1161 vdd a_n1358_n684# C3 w_n1316_n782# CMOSP w=7 l=3
+  ad=0 pd=0 as=0 ps=0
M1162 a_n844_n516# M gnd Gnd CMOSN w=5 l=2
+  ad=28 pd=22 as=0 ps=0
M1163 a_n797_n728# C1 a_n797_n761# Gnd CMOSN w=9 l=3
+  ad=72 pd=34 as=0 ps=0
M1164 vdd a_n2258_n792# a_n2045_n803# w_n2035_n704# CMOSP w=7 l=3
+  ad=0 pd=0 as=0 ps=0
M1165 a_n155_n657# M B0 w_n36_n486# CMOSP w=5 l=2
+  ad=60 pd=44 as=25 ps=20
M1166 a_n1358_n717# a_n1673_n776# gnd Gnd CMOSN w=9 l=3
+  ad=0 pd=0 as=0 ps=0
M1167 a_n155_n657# a_n44_n522# a_n15_n508# w_n36_n486# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1168 a_n955_n651# a_n844_n516# a_n815_n502# w_n836_n480# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1169 a_35_n684# M gnd Gnd CMOSN w=5 l=2
+  ad=28 pd=22 as=0 ps=0
M1170 a_n2472_n695# a_n2489_n709# a_n2460_n695# w_n2481_n673# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1171 a_n1515_n675# a_n1732_n679# gnd Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1172 C1 a_221_n679# a_278_n807# Gnd CMOSN w=9 l=3
+  ad=72 pd=34 as=0 ps=0
M1173 a_61_n771# a_3_n734# vdd vdd CMOSP w=5 l=3
+  ad=50 pd=30 as=0 ps=0
M1174 a_n894_n765# a_n952_n728# gnd Gnd CMOSN w=5 l=3
+  ad=40 pd=26 as=0 ps=0
M1175 a_n1720_n679# A2 vdd w_n1741_n657# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1176 a_n1732_n679# a_n1749_n693# A2 Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=23 ps=20
M1177 C1 a_274_n782# vdd w_263_n777# CMOSP w=7 l=3
+  ad=0 pd=0 as=0 ps=0
M1178 vdd a_n955_n651# a_n952_n728# w_n967_n731# CMOSP w=7 l=3
+  ad=0 pd=0 as=0 ps=0
M1179 a_n44_n522# M vdd w_n36_n486# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1180 a_n1673_n776# a_n1731_n739# vdd vdd CMOSP w=5 l=3
+  ad=50 pd=30 as=0 ps=0
M1181 a_n1749_n693# a_n1734_n662# gnd Gnd CMOSN w=5 l=2
+  ad=28 pd=22 as=0 ps=0
M1182 a_n579_n673# a_n894_n765# vdd w_n594_n676# CMOSP w=7 l=3
+  ad=0 pd=0 as=0 ps=0
M1183 a_n1301_n812# a_n1305_n787# gnd Gnd CMOSN w=9 l=3
+  ad=0 pd=0 as=0 ps=0
M1184 a_n1594_n513# B2 vdd w_n1615_n491# CMOSP w=5 l=2
+  ad=55 pd=42 as=0 ps=0
M1185 S3 a_n2284_n705# a_n2472_n695# Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1186 a_n526_n776# a_n739_n765# vdd w_n516_n677# CMOSP w=7 l=3
+  ad=0 pd=0 as=0 ps=0
M1187 a_n1734_n662# a_n1623_n527# a_n1594_n513# w_n1615_n491# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1188 S2 C2 a_n1732_n679# w_n1536_n653# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1189 a_221_n679# a_n94_n771# vdd w_206_n682# CMOSP w=7 l=3
+  ad=0 pd=0 as=0 ps=0
M1190 a_n2472_n695# a_n2474_n678# a_n2460_n695# Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1191 a_n1720_n679# A2 gnd Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
C0 w_n2355_n507# B3 10.81fF
C1 a_n1518_n776# vdd 1.53fF
C2 a_n2258_n792# vdd 1.53fF
C3 w_n2113_n703# vdd 2.26fF
C4 w_n2486_n758# vdd 2.26fF
C5 w_n1615_n491# a_n1623_n527# 4.79fF
C6 w_n836_n480# a_n844_n516# 4.79fF
C7 w_n2355_n507# a_n2363_n543# 4.79fF
C8 C2 gnd 0.90fF
C9 C3 gnd 0.90fF
C10 a_n2363_n543# B3 0.24fF
C11 w_n1746_n742# vdd 2.26fF
C12 w_n1373_n687# vdd 2.26fF
C13 w_n1615_n491# a_n1594_n513# 3.38fF
C14 a_35_n684# S0 0.24fF
C15 a_n953_n668# C1 0.36fF
C16 w_n812_n731# C1 2.66fF
C17 a_n2413_n792# vdd 0.99fF
C18 a_n1673_n776# vdd 0.99fF
C19 a_n1734_n662# gnd 0.58fF
C20 w_n2035_n704# vdd 2.26fF
C21 w_n757_n642# a_n736_n664# 3.38fF
C22 w_n1536_n653# S2 6.77fF
C23 w_n162_n652# a_n155_n657# 6.20fF
C24 w_n36_n486# B0 10.81fF
C25 w_n2481_n673# a_n2474_n678# 6.20fF
C26 w_n1615_n491# a_n1734_n662# 6.77fF
C27 C2 C1 0.72fF
C28 a_35_n684# a_n153_n674# 0.24fF
C29 w_n812_n731# a_n953_n668# 2.66fF
C30 w_n2276_n669# S3 6.77fF
C31 w_n836_n480# a_n815_n502# 3.38fF
C32 C1 S1 0.24fF
C33 w_n537_n771# a_n526_n776# 2.66fF
C34 w_n836_n480# a_n955_n651# 6.77fF
C35 C3 C2 0.72fF
C36 a_n1623_n527# a_n1734_n662# 0.39fF
C37 a_n955_n651# gnd 0.58fF
C38 M a_3_n734# 0.27fF
C39 w_n1591_n742# C2 2.66fF
C40 C1 a_221_n679# 0.27fF
C41 a_n739_n765# a_n526_n776# 0.27fF
C42 a_n1732_n679# C2 0.36fF
C43 w_n537_n771# a_n579_n673# 2.66fF
C44 a_n1734_n662# a_n1720_n679# 0.48fF
C45 a_n2472_n695# C3 0.36fF
C46 a_n44_n522# B0 0.24fF
C47 w_n1295_n688# a_n1305_n787# 0.56fF
C48 w_n2331_n758# C3 2.66fF
C49 a_n579_n673# a_n526_n776# 0.36fF
C50 a_n1518_n776# a_n1305_n787# 0.27fF
C51 a_n155_n657# a_n141_n674# 0.48fF
C52 a_n955_n651# a_n941_n668# 0.48fF
C53 a_n1734_n662# a_n1732_n679# 0.24fF
C54 w_n2056_n798# a_n2045_n803# 2.66fF
C55 w_n1591_n742# a_n1732_n679# 2.66fF
C56 a_n155_n657# a_n153_n674# 0.24fF
C57 a_n1358_n684# a_n1305_n787# 0.36fF
C58 C3 a_n1358_n684# 0.27fF
C59 a_n955_n651# a_n953_n668# 0.24fF
C60 a_n2284_n705# C3 0.15fF
C61 w_206_n682# a_221_n679# 0.56fF
C62 w_n2331_n758# a_n2472_n695# 2.66fF
C63 C2 a_n1673_n776# 0.54fF
C64 a_n765_n678# C1 0.15fF
C65 a_n2258_n792# a_n2045_n803# 0.27fF
C66 a_n2489_n709# a_n2472_n695# 0.24fF
C67 C3 a_n2413_n792# 0.54fF
C68 w_n2056_n798# a_n2098_n700# 2.66fF
C69 a_n844_n516# a_n955_n651# 0.39fF
C70 w_n1295_n688# a_n1518_n776# 5.32fF
C71 w_n1746_n742# a_n1734_n662# 2.66fF
C72 w_n967_n731# a_n955_n651# 2.66fF
C73 C2 a_n1515_n675# 0.48fF
C74 a_n2098_n700# a_n2045_n803# 0.36fF
C75 C3 a_n2255_n691# 0.48fF
C76 a_n1544_n689# C2 0.15fF
C77 a_n970_n682# a_n953_n668# 0.24fF
C78 a_n2284_n705# a_n2472_n695# 0.24fF
C79 a_n1734_n662# a_n1749_n693# 0.11fF
C80 a_n894_n765# a_n579_n673# 0.27fF
C81 a_n765_n678# a_n953_n668# 0.24fF
C82 a_n1749_n693# a_n1732_n679# 0.24fF
C83 w_n2035_n704# a_n2045_n803# 0.56fF
C84 w_n2113_n703# a_n2098_n700# 0.56fF
C85 a_n1732_n679# a_n1515_n675# 0.24fF
C86 a_n1544_n689# a_n1732_n679# 0.24fF
C87 a_n2472_n695# a_n2255_n691# 0.24fF
C88 w_n2035_n704# a_n2258_n792# 5.32fF
C89 w_n1373_n687# a_n1358_n684# 0.56fF
C90 w_n2113_n703# a_n2413_n792# 5.32fF
C91 a_n1673_n776# a_n1358_n684# 0.27fF
C92 a_n2413_n792# a_n2098_n700# 0.27fF
C93 w_n1373_n687# a_n1673_n776# 5.32fF
C94 a_n765_n678# S1 0.24fF
C95 w_43_n648# M 6.20fF
C96 w_284_n683# a_61_n771# 5.32fF
C97 w_n962_n646# A1 10.81fF
C98 a_3_n734# vdd 3.49fF
C99 a_n797_n728# vdd 3.49fF
C100 a_n2316_n755# vdd 3.49fF
C101 a_n952_n728# vdd 3.49fF
C102 a_n955_n651# a_n970_n682# 0.11fF
C103 S0 M 0.24fF
C104 w_n167_n737# A0 2.66fF
C105 a_n2471_n755# vdd 3.49fF
C106 a_n153_n674# M 0.36fF
C107 a_221_n679# a_274_n782# 0.36fF
C108 w_n2481_n673# A3 10.81fF
C109 a_n2334_n529# M 0.48fF
C110 C1 a_n797_n728# 0.27fF
C111 w_n12_n737# a_3_n734# 0.56fF
C112 a_n2474_n678# M 0.24fF
C113 w_n162_n652# vdd 3.38fF
C114 a_n170_n688# A0 0.24fF
C115 w_n757_n642# vdd 3.38fF
C116 a_n1720_n679# A2 0.24fF
C117 a_n1734_n662# A2 0.36fF
C118 a_n2474_n678# A3 0.36fF
C119 w_n812_n731# a_n797_n728# 0.56fF
C120 w_n962_n646# vdd 3.38fF
C121 a_n1732_n679# A2 0.72fF
C122 w_43_n648# vdd 3.38fF
C123 w_n1536_n653# vdd 3.38fF
C124 C3 a_n2316_n755# 0.27fF
C125 w_n967_n731# a_n952_n728# 0.56fF
C126 w_n1741_n657# vdd 3.38fF
C127 a_n15_n508# M 0.48fF
C128 w_n1746_n742# A2 2.66fF
C129 w_n2276_n669# vdd 3.38fF
C130 a_n155_n657# M 0.24fF
C131 a_n1749_n693# A2 0.24fF
C132 w_n2331_n758# a_n2316_n755# 0.56fF
C133 w_n2481_n673# vdd 3.38fF
C134 a_n155_n657# a_n152_n734# 0.27fF
C135 w_n757_n642# C1 6.20fF
C136 w_263_n777# vdd 2.26fF
C137 w_n2486_n758# a_n2471_n755# 0.56fF
C138 w_n537_n771# vdd 2.26fF
C139 a_n955_n651# a_n952_n728# 0.27fF
C140 w_n962_n646# a_n941_n668# 3.38fF
C141 w_n757_n642# a_n953_n668# 10.81fF
C142 w_n1316_n782# vdd 2.26fF
C143 w_n962_n646# a_n953_n668# 6.77fF
C144 w_43_n648# a_64_n670# 3.38fF
C145 a_n94_n771# vdd 0.99fF
C146 a_n739_n765# vdd 1.53fF
C147 w_284_n683# vdd 2.26fF
C148 w_n757_n642# S1 6.77fF
C149 w_n162_n652# a_n170_n688# 4.79fF
C150 w_n1536_n653# C2 6.20fF
C151 w_n1615_n491# B2 10.81fF
C152 w_263_n777# C1 0.56fF
C153 w_n12_n737# a_n153_n674# 2.66fF
C154 a_n894_n765# vdd 0.99fF
C155 a_n2474_n678# gnd 0.58fF
C156 w_n1741_n657# a_n1720_n679# 3.38fF
C157 w_n1536_n653# a_n1732_n679# 10.81fF
C158 w_n2276_n669# C3 6.20fF
C159 w_n1741_n657# a_n1734_n662# 6.20fF
C160 w_n2355_n507# a_n2334_n529# 3.38fF
C161 B3 a_n2334_n529# 0.24fF
C162 w_n1741_n657# a_n1732_n679# 6.77fF
C163 w_n836_n480# B1 10.81fF
C164 w_n2355_n507# a_n2474_n678# 6.77fF
C165 a_n153_n674# a_64_n670# 0.24fF
C166 B3 a_n2474_n678# 0.72fF
C167 a_n1623_n527# B2 0.24fF
C168 w_n2276_n669# a_n2472_n695# 10.81fF
C169 w_n2481_n673# a_n2460_n695# 3.38fF
C170 w_n962_n646# a_n955_n651# 6.20fF
C171 B2 a_n1594_n513# 0.24fF
C172 a_n2363_n543# a_n2474_n678# 0.39fF
C173 w_n36_n486# a_n15_n508# 3.38fF
C174 w_n2481_n673# a_n2472_n695# 6.77fF
C175 w_n537_n771# C2 0.56fF
C176 a_61_n771# vdd 1.53fF
C177 B2 a_n1734_n662# 0.72fF
C178 w_n1536_n653# a_n1515_n675# 3.38fF
C179 w_n2276_n669# a_n2284_n705# 4.79fF
C180 w_n757_n642# a_n765_n678# 4.79fF
C181 w_n962_n646# a_n970_n682# 4.79fF
C182 w_n1536_n653# a_n1544_n689# 4.79fF
C183 w_n1741_n657# a_n1749_n693# 4.79fF
C184 w_n2481_n673# a_n2489_n709# 4.79fF
C185 w_n36_n486# a_n155_n657# 6.77fF
C186 w_n516_n677# a_n526_n776# 0.56fF
C187 w_n1316_n782# a_n1305_n787# 2.66fF
C188 w_n1316_n782# C3 0.56fF
C189 a_n170_n688# a_n153_n674# 0.24fF
C190 C1 a_n894_n765# 0.54fF
C191 w_206_n682# a_n94_n771# 5.32fF
C192 a_n2474_n678# a_n2460_n695# 0.48fF
C193 a_n155_n657# gnd 0.58fF
C194 w_n2276_n669# a_n2255_n691# 3.38fF
C195 C1 a_n736_n664# 0.48fF
C196 a_n2474_n678# a_n2472_n695# 0.24fF
C197 w_n516_n677# a_n739_n765# 5.32fF
C198 a_n844_n516# B1 0.24fF
C199 C2 a_n579_n673# 0.27fF
C200 C2 S2 0.24fF
C201 w_263_n777# a_221_n679# 2.66fF
C202 C3 S3 0.24fF
C203 a_n2474_n678# a_n2489_n709# 0.11fF
C204 w_n2486_n758# a_n2474_n678# 2.66fF
C205 a_n953_n668# a_n736_n664# 0.24fF
C206 w_n594_n676# a_n579_n673# 0.56fF
C207 w_n1316_n782# a_n1358_n684# 2.66fF
C208 w_n167_n737# a_n155_n657# 2.66fF
C209 w_n594_n676# a_n894_n765# 5.32fF
C210 a_n44_n522# a_n155_n657# 0.39fF
C211 w_n162_n652# A0 10.81fF
C212 B1 a_n815_n502# 0.24fF
C213 a_n94_n771# a_221_n679# 0.27fF
C214 a_n2284_n705# S3 0.24fF
C215 B1 a_n955_n651# 0.72fF
C216 w_263_n777# a_274_n782# 2.66fF
C217 B0 a_n15_n508# 0.24fF
C218 a_n155_n657# a_n170_n688# 0.11fF
C219 a_n152_n734# vdd 3.49fF
C220 a_n1544_n689# S2 0.24fF
C221 B0 a_n155_n657# 0.72fF
C222 w_n36_n486# M 6.20fF
C223 a_n1576_n739# vdd 3.49fF
C224 w_n836_n480# M 6.20fF
C225 a_n141_n674# A0 0.24fF
C226 a_n1731_n739# vdd 3.49fF
C227 w_284_n683# a_274_n782# 0.56fF
C228 w_n1615_n491# M 6.20fF
C229 w_n1741_n657# A2 10.81fF
C230 a_n153_n674# A0 0.72fF
C231 w_n2355_n507# M 6.20fF
C232 w_n12_n737# M 2.66fF
C233 a_64_n670# M 0.48fF
C234 a_n941_n668# A1 0.24fF
C235 w_n167_n737# a_n152_n734# 0.56fF
C236 a_n953_n668# A1 0.72fF
C237 a_n1594_n513# M 0.48fF
C238 a_61_n771# a_274_n782# 0.27fF
C239 a_n1734_n662# M 0.24fF
C240 w_n967_n731# A1 2.66fF
C241 C2 a_n1576_n739# 0.27fF
C242 a_n2460_n695# A3 0.24fF
C243 w_n36_n486# vdd 3.38fF
C244 a_n2472_n695# A3 0.72fF
C245 a_n155_n657# A0 0.36fF
C246 a_n815_n502# M 0.48fF
C247 w_n1591_n742# a_n1576_n739# 0.56fF
C248 w_n836_n480# vdd 3.38fF
C249 a_n955_n651# M 0.24fF
C250 a_n2489_n709# A3 0.24fF
C251 w_n2056_n798# carry 0.56fF
C252 a_n2474_n678# a_n2471_n755# 0.27fF
C253 a_n1734_n662# a_n1731_n739# 0.27fF
C254 w_n2486_n758# A3 2.66fF
C255 w_n1615_n491# vdd 3.38fF
C256 a_n955_n651# A1 0.36fF
C257 w_n162_n652# a_n141_n674# 3.38fF
C258 w_n2355_n507# vdd 3.38fF
C259 w_n12_n737# vdd 2.26fF
C260 w_n162_n652# a_n153_n674# 6.77fF
C261 w_43_n648# S0 6.77fF
C262 a_n2098_n700# carry 0.27fF
C263 a_n970_n682# A1 0.24fF
C264 w_n167_n737# vdd 2.26fF
C265 w_n1746_n742# a_n1731_n739# 0.56fF
C266 w_206_n682# vdd 2.26fF
C267 w_n812_n731# vdd 2.26fF
C268 w_43_n648# a_n153_n674# 10.81fF
C269 w_n967_n731# vdd 2.26fF
C270 w_n516_n677# vdd 2.26fF
C271 C1 gnd 0.90fF
C272 w_n2056_n798# vdd 2.26fF
C273 w_n1591_n742# vdd 2.26fF
C274 w_n594_n676# vdd 2.26fF
C275 w_n36_n486# a_n44_n522# 4.79fF
C276 w_43_n648# a_35_n684# 4.79fF
C277 w_n2331_n758# vdd 2.26fF
C278 w_n1295_n688# vdd 2.26fF
C279 gnd Gnd 225.37fF
C280 vdd Gnd 265.83fF
C281 carry Gnd 7.29fF
C282 a_3_n734# Gnd 7.47fF
C283 M Gnd 157.36fF
C284 a_n152_n734# Gnd 7.10fF
C285 A0 Gnd 33.52fF
C286 a_n2316_n755# Gnd 21.61fF
C287 a_n2471_n755# Gnd 1.32fF
C288 A3 Gnd 34.27fF
C289 a_n1576_n739# Gnd 21.61fF
C290 a_n1731_n739# Gnd 21.61fF
C291 A2 Gnd 34.27fF
C292 a_n797_n728# Gnd 21.61fF
C293 a_n952_n728# Gnd 7.10fF
C294 A1 Gnd 33.70fF
C295 a_274_n782# Gnd 41.71fF
C296 a_61_n771# Gnd 46.16fF
C297 a_221_n679# Gnd 34.24fF
C298 a_n94_n771# Gnd 90.05fF
C299 a_64_n670# Gnd 15.09fF
C300 S0 Gnd 12.69fF
C301 a_n141_n674# Gnd 15.09fF
C302 a_n153_n674# Gnd 73.29fF
C303 a_n526_n776# Gnd 41.71fF
C304 a_n739_n765# Gnd 46.16fF
C305 a_n579_n673# Gnd 34.24fF
C306 a_n894_n765# Gnd 90.05fF
C307 a_n736_n664# Gnd 15.09fF
C308 S1 Gnd 12.69fF
C309 a_n170_n688# Gnd 71.09fF
C310 a_35_n684# Gnd 71.09fF
C311 C1 Gnd 269.74fF
C312 a_n941_n668# Gnd 15.09fF
C313 a_n953_n668# Gnd 73.29fF
C314 a_n1305_n787# Gnd 41.71fF
C315 a_n2045_n803# Gnd 41.71fF
C316 a_n1518_n776# Gnd 46.16fF
C317 a_n1358_n684# Gnd 34.24fF
C318 a_n1673_n776# Gnd 90.05fF
C319 a_n1515_n675# Gnd 15.09fF
C320 S2 Gnd 12.69fF
C321 C2 Gnd 414.84fF
C322 a_n1720_n679# Gnd 15.09fF
C323 a_n1732_n679# Gnd 73.29fF
C324 a_n2258_n792# Gnd 46.16fF
C325 a_n2098_n700# Gnd 34.24fF
C326 a_n2413_n792# Gnd 90.05fF
C327 a_n2255_n691# Gnd 15.09fF
C328 S3 Gnd 12.69fF
C329 C3 Gnd 411.95fF
C330 a_n2460_n695# Gnd 15.09fF
C331 a_n2472_n695# Gnd 73.29fF
C332 a_n2489_n709# Gnd 71.09fF
C333 a_n2284_n705# Gnd 19.36fF
C334 a_n1749_n693# Gnd 71.09fF
C335 a_n1544_n689# Gnd 71.09fF
C336 a_n970_n682# Gnd 71.09fF
C337 a_n765_n678# Gnd 71.09fF
C338 a_n15_n508# Gnd 15.09fF
C339 a_n155_n657# Gnd 101.01fF
C340 B0 Gnd 24.28fF
C341 a_n815_n502# Gnd 15.09fF
C342 a_n955_n651# Gnd 101.01fF
C343 B1 Gnd 24.28fF
C344 a_n44_n522# Gnd 71.09fF
C345 a_n1594_n513# Gnd 15.09fF
C346 a_n1734_n662# Gnd 101.01fF
C347 B2 Gnd 24.28fF
C348 a_n2334_n529# Gnd 15.09fF
C349 a_n2474_n678# Gnd 101.01fF
C350 B3 Gnd 24.28fF
C351 a_n2363_n543# Gnd 71.09fF
C352 a_n1623_n527# Gnd 71.09fF
C353 a_n844_n516# Gnd 71.09fF

.tran 0.1n 800n

.control
run 

*  plot v(B0)+4 v(M)+2 
* plot v(out)
* plot v(B0)+6 v(A0)+4 v(C1)+2 v(S0)  
* plot v(B1)+8 v(A1)+6 v(C1)+4 v(C2)+2 v(S1)  

plot v(carry)+8 v(S3)+6 v(S2)+4 v(S1)+2 v(S0)
* plot v(C3)+4 v(C2)+2 v(C1)
* plot v(A1)+2 v(A0)
* plot v(xor_check)+6 v(A0)+4 v(M)+2 v(C1)  


.endc

.end
