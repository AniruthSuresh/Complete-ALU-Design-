magic
tech scmos
timestamp 1699736150
<< nwell >>
rect 238 137 276 153
rect 290 135 331 153
rect 133 41 174 59
rect 240 54 278 70
rect 292 52 333 70
rect 134 -56 175 -38
rect 238 -46 276 -30
rect 290 -48 331 -30
rect 239 -135 277 -119
rect 291 -137 332 -119
<< polysilicon >>
rect 250 147 253 151
rect 261 147 264 151
rect 308 147 311 150
rect 250 136 253 140
rect 250 116 253 132
rect 261 128 264 140
rect 308 127 311 142
rect 261 116 264 124
rect 308 108 311 123
rect 250 104 253 107
rect 261 104 264 107
rect 308 99 311 103
rect 252 64 255 68
rect 263 64 266 68
rect 310 64 313 67
rect 151 53 154 56
rect 252 53 255 57
rect 151 33 154 48
rect 252 33 255 49
rect 263 45 266 57
rect 310 44 313 59
rect 263 33 266 41
rect 151 14 154 29
rect 310 25 313 40
rect 252 21 255 24
rect 263 21 266 24
rect 310 16 313 20
rect 151 5 154 9
rect 250 -36 253 -32
rect 261 -36 264 -32
rect 308 -36 311 -33
rect 152 -44 155 -41
rect 250 -47 253 -43
rect 152 -64 155 -49
rect 250 -67 253 -51
rect 261 -55 264 -43
rect 308 -56 311 -41
rect 261 -67 264 -59
rect 152 -83 155 -68
rect 308 -75 311 -60
rect 250 -79 253 -76
rect 261 -79 264 -76
rect 308 -84 311 -80
rect 152 -92 155 -88
rect 251 -125 254 -121
rect 262 -125 265 -121
rect 309 -125 312 -122
rect 251 -136 254 -132
rect 251 -156 254 -140
rect 262 -144 265 -132
rect 309 -145 312 -130
rect 262 -156 265 -148
rect 309 -164 312 -149
rect 251 -168 254 -165
rect 262 -168 265 -165
rect 309 -173 312 -169
<< ndiffusion >>
rect 248 112 250 116
rect 244 107 250 112
rect 253 107 261 116
rect 264 112 267 116
rect 271 112 272 116
rect 264 107 272 112
rect 305 103 308 108
rect 311 103 315 108
rect 250 29 252 33
rect 246 24 252 29
rect 255 24 263 33
rect 266 29 269 33
rect 273 29 274 33
rect 266 24 274 29
rect 307 20 310 25
rect 313 20 317 25
rect 148 9 151 14
rect 154 9 158 14
rect 248 -71 250 -67
rect 244 -76 250 -71
rect 253 -76 261 -67
rect 264 -71 267 -67
rect 271 -71 272 -67
rect 264 -76 272 -71
rect 305 -80 308 -75
rect 311 -80 315 -75
rect 149 -88 152 -83
rect 155 -88 159 -83
rect 249 -160 251 -156
rect 245 -165 251 -160
rect 254 -165 262 -156
rect 265 -160 268 -156
rect 272 -160 273 -156
rect 265 -165 273 -160
rect 306 -169 309 -164
rect 312 -169 316 -164
<< pdiffusion >>
rect 247 143 250 147
rect 243 140 250 143
rect 253 143 256 147
rect 260 143 261 147
rect 253 140 261 143
rect 264 143 267 147
rect 264 140 271 143
rect 304 142 308 147
rect 311 142 315 147
rect 319 142 321 147
rect 249 60 252 64
rect 245 57 252 60
rect 255 60 258 64
rect 262 60 263 64
rect 255 57 263 60
rect 266 60 269 64
rect 266 57 273 60
rect 306 59 310 64
rect 313 59 317 64
rect 321 59 323 64
rect 147 48 151 53
rect 154 48 158 53
rect 162 48 164 53
rect 247 -40 250 -36
rect 243 -43 250 -40
rect 253 -40 256 -36
rect 260 -40 261 -36
rect 253 -43 261 -40
rect 264 -40 267 -36
rect 264 -43 271 -40
rect 304 -41 308 -36
rect 311 -41 315 -36
rect 319 -41 321 -36
rect 148 -49 152 -44
rect 155 -49 159 -44
rect 163 -49 165 -44
rect 248 -129 251 -125
rect 244 -132 251 -129
rect 254 -129 257 -125
rect 261 -129 262 -125
rect 254 -132 262 -129
rect 265 -129 268 -125
rect 265 -132 272 -129
rect 305 -130 309 -125
rect 312 -130 316 -125
rect 320 -130 322 -125
<< metal1 >>
rect 243 153 303 157
rect 307 153 332 157
rect 243 147 247 153
rect 267 147 271 153
rect 300 147 303 153
rect 256 136 260 143
rect 204 132 249 136
rect 256 133 271 136
rect 133 59 146 63
rect 150 59 174 63
rect 143 53 146 59
rect 130 29 150 33
rect 159 31 162 48
rect 204 31 208 132
rect 267 130 271 133
rect 159 26 208 31
rect 159 14 162 26
rect 143 2 147 9
rect 133 -4 175 2
rect 134 -38 147 -34
rect 151 -38 175 -34
rect 144 -44 147 -38
rect 160 -64 163 -49
rect 204 -47 208 26
rect 224 124 260 128
rect 267 127 272 130
rect 224 45 228 124
rect 267 123 307 127
rect 267 116 271 123
rect 244 103 248 112
rect 316 108 319 142
rect 244 101 290 103
rect 300 101 304 103
rect 244 100 304 101
rect 272 98 304 100
rect 245 70 305 74
rect 309 70 334 74
rect 245 64 249 70
rect 269 64 273 70
rect 302 64 305 70
rect 258 53 262 60
rect 243 49 251 53
rect 258 50 273 53
rect 269 47 273 50
rect 224 41 262 45
rect 269 44 274 47
rect 204 -51 206 -47
rect 224 -64 228 41
rect 269 40 309 44
rect 269 33 273 40
rect 246 20 250 29
rect 318 25 321 59
rect 246 17 292 20
rect 274 16 292 17
rect 302 16 306 20
rect 274 12 306 16
rect 243 -30 303 -26
rect 307 -30 332 -26
rect 243 -36 247 -30
rect 267 -36 271 -30
rect 300 -36 303 -30
rect 256 -47 260 -40
rect 243 -51 249 -47
rect 256 -50 271 -47
rect 267 -53 271 -50
rect 119 -68 151 -64
rect 160 -67 228 -64
rect 233 -59 260 -55
rect 267 -56 272 -53
rect 119 -110 123 -68
rect 160 -83 163 -67
rect 144 -95 148 -88
rect 134 -101 176 -95
rect 233 -110 237 -59
rect 267 -60 307 -56
rect 267 -67 271 -60
rect 244 -80 248 -71
rect 316 -75 319 -41
rect 244 -82 290 -80
rect 300 -82 304 -80
rect 244 -83 304 -82
rect 272 -85 304 -83
rect 119 -114 237 -110
rect 217 -144 221 -114
rect 244 -119 304 -115
rect 308 -119 333 -115
rect 244 -125 248 -119
rect 268 -125 272 -119
rect 301 -125 304 -119
rect 257 -136 261 -129
rect 244 -140 250 -136
rect 257 -139 272 -136
rect 268 -142 272 -139
rect 217 -148 261 -144
rect 268 -145 273 -142
rect 268 -149 308 -145
rect 268 -156 272 -149
rect 245 -169 249 -160
rect 317 -164 320 -130
rect 245 -171 291 -169
rect 301 -171 305 -169
rect 245 -172 305 -171
rect 273 -175 305 -172
<< metal2 >>
rect 126 68 234 72
rect 126 49 130 68
rect 230 53 234 68
rect 230 49 239 53
rect 99 45 130 49
rect 99 -136 103 45
rect 126 33 130 45
rect 211 -51 238 -47
rect 99 -140 240 -136
<< ntransistor >>
rect 250 107 253 116
rect 261 107 264 116
rect 308 103 311 108
rect 252 24 255 33
rect 263 24 266 33
rect 310 20 313 25
rect 151 9 154 14
rect 250 -76 253 -67
rect 261 -76 264 -67
rect 308 -80 311 -75
rect 152 -88 155 -83
rect 251 -165 254 -156
rect 262 -165 265 -156
rect 309 -169 312 -164
<< ptransistor >>
rect 250 140 253 147
rect 261 140 264 147
rect 308 142 311 147
rect 252 57 255 64
rect 263 57 266 64
rect 310 59 313 64
rect 151 48 154 53
rect 250 -43 253 -36
rect 261 -43 264 -36
rect 308 -41 311 -36
rect 152 -49 155 -44
rect 251 -132 254 -125
rect 262 -132 265 -125
rect 309 -130 312 -125
<< polycontact >>
rect 249 132 253 136
rect 260 124 264 128
rect 307 123 311 127
rect 251 49 255 53
rect 262 41 266 45
rect 309 40 313 44
rect 150 29 154 33
rect 249 -51 253 -47
rect 151 -68 155 -64
rect 260 -59 264 -55
rect 307 -60 311 -56
rect 250 -140 254 -136
rect 261 -148 265 -144
rect 308 -149 312 -145
<< ndcontact >>
rect 244 112 248 116
rect 267 112 271 116
rect 300 103 305 108
rect 315 103 319 108
rect 246 29 250 33
rect 269 29 273 33
rect 302 20 307 25
rect 317 20 321 25
rect 143 9 148 14
rect 158 9 162 14
rect 244 -71 248 -67
rect 267 -71 271 -67
rect 300 -80 305 -75
rect 315 -80 319 -75
rect 144 -88 149 -83
rect 159 -88 163 -83
rect 245 -160 249 -156
rect 268 -160 272 -156
rect 301 -169 306 -164
rect 316 -169 320 -164
<< pdcontact >>
rect 243 143 247 147
rect 256 143 260 147
rect 267 143 271 147
rect 300 142 304 147
rect 315 142 319 147
rect 245 60 249 64
rect 258 60 262 64
rect 269 60 273 64
rect 302 59 306 64
rect 317 59 321 64
rect 143 48 147 53
rect 158 48 162 53
rect 243 -40 247 -36
rect 256 -40 260 -36
rect 267 -40 271 -36
rect 300 -41 304 -36
rect 315 -41 319 -36
rect 144 -49 148 -44
rect 159 -49 163 -44
rect 244 -129 248 -125
rect 257 -129 261 -125
rect 268 -129 272 -125
rect 301 -130 305 -125
rect 316 -130 320 -125
<< m2contact >>
rect 126 29 130 33
rect 239 49 243 53
rect 206 -51 211 -47
rect 238 -51 243 -47
rect 240 -140 244 -136
<< nsubstratencontact >>
rect 303 153 307 157
rect 305 70 309 74
rect 146 59 150 63
rect 303 -30 307 -26
rect 147 -38 151 -34
rect 304 -119 308 -115
<< labels >>
rlabel metal1 156 61 156 61 5 vdd
rlabel metal1 151 -1 151 -1 1 gnd
rlabel metal1 157 -36 157 -36 5 vdd
rlabel metal1 152 -98 152 -98 1 gnd
rlabel metal1 144 31 144 31 1 A0
rlabel metal1 145 -65 145 -65 1 A1
rlabel metal1 286 72 286 72 1 vdd
rlabel metal1 282 -28 282 -28 1 vdd
rlabel metal1 283 -116 283 -116 1 vdd
rlabel metal1 286 -172 286 -172 1 gnd
rlabel metal1 281 -83 281 -83 1 gnd
rlabel metal1 280 15 280 15 1 gnd
rlabel metal1 284 100 284 100 1 gnd
rlabel metal1 317 126 317 126 1 D0
rlabel metal1 319 42 319 42 1 D1
rlabel metal1 318 -58 318 -58 1 D2
rlabel metal1 318 -149 318 -149 1 D3
rlabel metal1 282 155 282 155 5 vdd
<< end >>
