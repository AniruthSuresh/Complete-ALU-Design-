magic
tech scmos
timestamp 1699729768
<< nwell >>
rect -2355 -507 -2275 -484
rect -1615 -491 -1535 -468
rect -836 -480 -756 -457
rect -156 -486 -76 -463
rect -2481 -673 -2401 -650
rect -2276 -669 -2196 -646
rect -1741 -657 -1661 -634
rect -1536 -653 -1456 -630
rect -962 -646 -882 -623
rect -757 -642 -677 -619
rect -282 -652 -202 -629
rect -77 -648 3 -625
rect -1373 -687 -1335 -671
rect -2113 -703 -2075 -687
rect -1295 -688 -1257 -672
rect -594 -676 -556 -660
rect -516 -677 -478 -661
rect 86 -682 124 -666
rect 164 -683 202 -667
rect -2035 -704 -1997 -688
rect -1746 -742 -1708 -726
rect -2486 -758 -2448 -742
rect -2434 -760 -2393 -742
rect -2331 -758 -2293 -742
rect -2279 -760 -2238 -742
rect -1694 -744 -1653 -726
rect -1591 -742 -1553 -726
rect -1539 -744 -1498 -726
rect -967 -731 -929 -715
rect -915 -733 -874 -715
rect -812 -731 -774 -715
rect -760 -733 -719 -715
rect -287 -737 -249 -721
rect -235 -739 -194 -721
rect -132 -737 -94 -721
rect -80 -739 -39 -721
rect -1316 -782 -1278 -766
rect -537 -771 -499 -755
rect 143 -777 181 -761
rect -2056 -798 -2018 -782
<< polysilicon >>
rect -844 -437 -808 -435
rect -1623 -448 -1587 -446
rect -2363 -464 -2327 -462
rect -2363 -541 -2361 -464
rect -2348 -493 -2346 -491
rect -2329 -493 -2327 -464
rect -2304 -493 -2302 -491
rect -2285 -493 -2283 -491
rect -2348 -510 -2346 -498
rect -2329 -500 -2327 -498
rect -2304 -510 -2302 -498
rect -2285 -510 -2283 -498
rect -2348 -512 -2327 -510
rect -2348 -524 -2346 -521
rect -2329 -524 -2327 -512
rect -2303 -514 -2302 -510
rect -2284 -514 -2283 -510
rect -2274 -513 -2268 -511
rect -2304 -524 -2302 -514
rect -2285 -524 -2283 -514
rect -2348 -541 -2346 -529
rect -2329 -537 -2327 -529
rect -2304 -531 -2302 -529
rect -2285 -537 -2283 -529
rect -2329 -539 -2283 -537
rect -2270 -541 -2268 -513
rect -1623 -525 -1621 -448
rect -1608 -477 -1606 -475
rect -1589 -477 -1587 -448
rect -1564 -477 -1562 -475
rect -1545 -477 -1543 -475
rect -1608 -494 -1606 -482
rect -1589 -484 -1587 -482
rect -1564 -494 -1562 -482
rect -1545 -494 -1543 -482
rect -1608 -496 -1587 -494
rect -1608 -508 -1606 -505
rect -1589 -508 -1587 -496
rect -1563 -498 -1562 -494
rect -1544 -498 -1543 -494
rect -1534 -497 -1528 -495
rect -1564 -508 -1562 -498
rect -1545 -508 -1543 -498
rect -1608 -525 -1606 -513
rect -1589 -521 -1587 -513
rect -1564 -515 -1562 -513
rect -1545 -521 -1543 -513
rect -1589 -523 -1543 -521
rect -1530 -525 -1528 -497
rect -844 -514 -842 -437
rect -829 -466 -827 -464
rect -810 -466 -808 -437
rect -164 -443 -128 -441
rect -785 -466 -783 -464
rect -766 -466 -764 -464
rect -829 -483 -827 -471
rect -810 -473 -808 -471
rect -785 -483 -783 -471
rect -766 -483 -764 -471
rect -829 -485 -808 -483
rect -829 -497 -827 -494
rect -810 -497 -808 -485
rect -784 -487 -783 -483
rect -765 -487 -764 -483
rect -755 -486 -749 -484
rect -785 -497 -783 -487
rect -766 -497 -764 -487
rect -829 -514 -827 -502
rect -810 -510 -808 -502
rect -785 -504 -783 -502
rect -766 -510 -764 -502
rect -810 -512 -764 -510
rect -751 -514 -749 -486
rect -844 -516 -749 -514
rect -164 -520 -162 -443
rect -149 -472 -147 -470
rect -130 -472 -128 -443
rect -105 -472 -103 -470
rect -86 -472 -84 -470
rect -149 -489 -147 -477
rect -130 -479 -128 -477
rect -105 -489 -103 -477
rect -86 -489 -84 -477
rect -149 -491 -128 -489
rect -149 -503 -147 -500
rect -130 -503 -128 -491
rect -104 -493 -103 -489
rect -85 -493 -84 -489
rect -75 -492 -69 -490
rect -105 -503 -103 -493
rect -86 -503 -84 -493
rect -149 -520 -147 -508
rect -130 -516 -128 -508
rect -105 -510 -103 -508
rect -86 -516 -84 -508
rect -130 -518 -84 -516
rect -71 -520 -69 -492
rect -164 -522 -69 -520
rect -1623 -527 -1528 -525
rect -2363 -543 -2268 -541
rect -765 -599 -729 -597
rect -970 -603 -934 -601
rect -1544 -610 -1508 -608
rect -1749 -614 -1713 -612
rect -2284 -626 -2248 -624
rect -2489 -630 -2453 -628
rect -2489 -707 -2487 -630
rect -2474 -659 -2472 -657
rect -2455 -659 -2453 -630
rect -2430 -659 -2428 -657
rect -2411 -659 -2409 -657
rect -2474 -676 -2472 -664
rect -2455 -666 -2453 -664
rect -2430 -676 -2428 -664
rect -2474 -678 -2453 -676
rect -2474 -690 -2472 -687
rect -2455 -690 -2453 -678
rect -2429 -680 -2428 -676
rect -2411 -677 -2409 -664
rect -2430 -690 -2428 -680
rect -2410 -681 -2409 -677
rect -2400 -679 -2394 -677
rect -2411 -690 -2409 -681
rect -2474 -707 -2472 -695
rect -2455 -703 -2453 -695
rect -2430 -697 -2428 -695
rect -2411 -703 -2409 -695
rect -2455 -705 -2409 -703
rect -2396 -707 -2394 -679
rect -2284 -703 -2282 -626
rect -2269 -655 -2267 -653
rect -2250 -655 -2248 -626
rect -2225 -655 -2223 -653
rect -2206 -655 -2204 -653
rect -2269 -672 -2267 -660
rect -2250 -662 -2248 -660
rect -2225 -672 -2223 -660
rect -2206 -672 -2204 -660
rect -2269 -674 -2248 -672
rect -2269 -686 -2267 -683
rect -2250 -686 -2248 -674
rect -2224 -676 -2223 -672
rect -2205 -676 -2204 -672
rect -2195 -675 -2189 -673
rect -2225 -686 -2223 -676
rect -2206 -686 -2204 -676
rect -2269 -703 -2267 -691
rect -2250 -699 -2248 -691
rect -2225 -693 -2223 -691
rect -2206 -699 -2204 -691
rect -2250 -701 -2204 -699
rect -2191 -703 -2189 -675
rect -2101 -693 -2098 -689
rect -2090 -693 -2087 -689
rect -2023 -694 -2020 -690
rect -2012 -694 -2009 -690
rect -1749 -691 -1747 -614
rect -1734 -643 -1732 -641
rect -1715 -643 -1713 -614
rect -1690 -643 -1688 -641
rect -1671 -643 -1669 -641
rect -1734 -660 -1732 -648
rect -1715 -650 -1713 -648
rect -1690 -660 -1688 -648
rect -1734 -662 -1713 -660
rect -1734 -674 -1732 -671
rect -1715 -674 -1713 -662
rect -1689 -664 -1688 -660
rect -1671 -661 -1669 -648
rect -1690 -674 -1688 -664
rect -1670 -665 -1669 -661
rect -1660 -663 -1654 -661
rect -1671 -674 -1669 -665
rect -1734 -691 -1732 -679
rect -1715 -687 -1713 -679
rect -1690 -681 -1688 -679
rect -1671 -687 -1669 -679
rect -1715 -689 -1669 -687
rect -1656 -691 -1654 -663
rect -1544 -687 -1542 -610
rect -1529 -639 -1527 -637
rect -1510 -639 -1508 -610
rect -1485 -639 -1483 -637
rect -1466 -639 -1464 -637
rect -1529 -656 -1527 -644
rect -1510 -646 -1508 -644
rect -1485 -656 -1483 -644
rect -1466 -656 -1464 -644
rect -1529 -658 -1508 -656
rect -1529 -670 -1527 -667
rect -1510 -670 -1508 -658
rect -1484 -660 -1483 -656
rect -1465 -660 -1464 -656
rect -1455 -659 -1449 -657
rect -1485 -670 -1483 -660
rect -1466 -670 -1464 -660
rect -1529 -687 -1527 -675
rect -1510 -683 -1508 -675
rect -1485 -677 -1483 -675
rect -1466 -683 -1464 -675
rect -1510 -685 -1464 -683
rect -1451 -687 -1449 -659
rect -1361 -677 -1358 -673
rect -1350 -677 -1347 -673
rect -1283 -678 -1280 -674
rect -1272 -678 -1269 -674
rect -1544 -689 -1449 -687
rect -1361 -688 -1358 -684
rect -1749 -693 -1654 -691
rect -2284 -705 -2189 -703
rect -2101 -704 -2098 -700
rect -2489 -709 -2394 -707
rect -2101 -724 -2098 -708
rect -2090 -712 -2087 -700
rect -2023 -705 -2020 -701
rect -2090 -724 -2087 -716
rect -2023 -725 -2020 -709
rect -2012 -713 -2009 -701
rect -1361 -708 -1358 -692
rect -1350 -696 -1347 -684
rect -970 -680 -968 -603
rect -955 -632 -953 -630
rect -936 -632 -934 -603
rect -911 -632 -909 -630
rect -892 -632 -890 -630
rect -955 -649 -953 -637
rect -936 -639 -934 -637
rect -911 -649 -909 -637
rect -955 -651 -934 -649
rect -955 -663 -953 -660
rect -936 -663 -934 -651
rect -910 -653 -909 -649
rect -892 -650 -890 -637
rect -911 -663 -909 -653
rect -891 -654 -890 -650
rect -881 -652 -875 -650
rect -892 -663 -890 -654
rect -955 -680 -953 -668
rect -936 -676 -934 -668
rect -911 -670 -909 -668
rect -892 -676 -890 -668
rect -936 -678 -890 -676
rect -877 -680 -875 -652
rect -765 -676 -763 -599
rect -750 -628 -748 -626
rect -731 -628 -729 -599
rect -85 -605 -49 -603
rect -290 -609 -254 -607
rect -706 -628 -704 -626
rect -687 -628 -685 -626
rect -750 -645 -748 -633
rect -731 -635 -729 -633
rect -706 -645 -704 -633
rect -687 -645 -685 -633
rect -750 -647 -729 -645
rect -750 -659 -748 -656
rect -731 -659 -729 -647
rect -705 -649 -704 -645
rect -686 -649 -685 -645
rect -676 -648 -670 -646
rect -706 -659 -704 -649
rect -687 -659 -685 -649
rect -750 -676 -748 -664
rect -731 -672 -729 -664
rect -706 -666 -704 -664
rect -687 -672 -685 -664
rect -731 -674 -685 -672
rect -672 -676 -670 -648
rect -582 -666 -579 -662
rect -571 -666 -568 -662
rect -504 -667 -501 -663
rect -493 -667 -490 -663
rect -765 -678 -670 -676
rect -582 -677 -579 -673
rect -970 -682 -875 -680
rect -1283 -689 -1280 -685
rect -1350 -708 -1347 -700
rect -1283 -709 -1280 -693
rect -1272 -697 -1269 -685
rect -582 -697 -579 -681
rect -571 -685 -568 -673
rect -504 -678 -501 -674
rect -571 -697 -568 -689
rect -1272 -709 -1269 -701
rect -504 -698 -501 -682
rect -493 -686 -490 -674
rect -290 -686 -288 -609
rect -275 -638 -273 -636
rect -256 -638 -254 -609
rect -231 -638 -229 -636
rect -212 -638 -210 -636
rect -275 -655 -273 -643
rect -256 -645 -254 -643
rect -231 -655 -229 -643
rect -275 -657 -254 -655
rect -275 -669 -273 -666
rect -256 -669 -254 -657
rect -230 -659 -229 -655
rect -212 -656 -210 -643
rect -231 -669 -229 -659
rect -211 -660 -210 -656
rect -201 -658 -195 -656
rect -212 -669 -210 -660
rect -275 -686 -273 -674
rect -256 -682 -254 -674
rect -231 -676 -229 -674
rect -212 -682 -210 -674
rect -256 -684 -210 -682
rect -197 -686 -195 -658
rect -85 -682 -83 -605
rect -70 -634 -68 -632
rect -51 -634 -49 -605
rect -26 -634 -24 -632
rect -7 -634 -5 -632
rect -70 -651 -68 -639
rect -51 -641 -49 -639
rect -26 -651 -24 -639
rect -7 -651 -5 -639
rect -70 -653 -49 -651
rect -70 -665 -68 -662
rect -51 -665 -49 -653
rect -25 -655 -24 -651
rect -6 -655 -5 -651
rect 4 -654 10 -652
rect -26 -665 -24 -655
rect -7 -665 -5 -655
rect -70 -682 -68 -670
rect -51 -678 -49 -670
rect -26 -672 -24 -670
rect -7 -678 -5 -670
rect -51 -680 -5 -678
rect 8 -682 10 -654
rect 98 -672 101 -668
rect 109 -672 112 -668
rect 176 -673 179 -669
rect 187 -673 190 -669
rect -85 -684 10 -682
rect 98 -683 101 -679
rect -290 -688 -195 -686
rect -493 -698 -490 -690
rect -582 -709 -579 -706
rect -571 -709 -568 -706
rect 98 -703 101 -687
rect 109 -691 112 -679
rect 176 -684 179 -680
rect 109 -703 112 -695
rect -2012 -725 -2009 -717
rect -1361 -720 -1358 -717
rect -1350 -720 -1347 -717
rect -504 -710 -501 -707
rect -493 -710 -490 -707
rect 176 -704 179 -688
rect 187 -692 190 -680
rect 187 -704 190 -696
rect 98 -715 101 -712
rect 109 -715 112 -712
rect 176 -716 179 -713
rect 187 -716 190 -713
rect -1283 -721 -1280 -718
rect -1272 -721 -1269 -718
rect -955 -721 -952 -717
rect -944 -721 -941 -717
rect -897 -721 -894 -718
rect -800 -721 -797 -717
rect -789 -721 -786 -717
rect -742 -721 -739 -718
rect -2101 -736 -2098 -733
rect -2090 -736 -2087 -733
rect -1734 -732 -1731 -728
rect -1723 -732 -1720 -728
rect -1676 -732 -1673 -729
rect -1579 -732 -1576 -728
rect -1568 -732 -1565 -728
rect -1521 -732 -1518 -729
rect -955 -732 -952 -728
rect -2023 -737 -2020 -734
rect -2012 -737 -2009 -734
rect -1734 -743 -1731 -739
rect -2474 -748 -2471 -744
rect -2463 -748 -2460 -744
rect -2416 -748 -2413 -745
rect -2319 -748 -2316 -744
rect -2308 -748 -2305 -744
rect -2261 -748 -2258 -745
rect -2474 -759 -2471 -755
rect -2474 -779 -2471 -763
rect -2463 -767 -2460 -755
rect -2416 -768 -2413 -753
rect -2319 -759 -2316 -755
rect -2463 -779 -2460 -771
rect -2416 -787 -2413 -772
rect -2319 -779 -2316 -763
rect -2308 -767 -2305 -755
rect -2261 -768 -2258 -753
rect -1734 -763 -1731 -747
rect -1723 -751 -1720 -739
rect -1676 -752 -1673 -737
rect -1579 -743 -1576 -739
rect -1723 -763 -1720 -755
rect -2308 -779 -2305 -771
rect -1676 -771 -1673 -756
rect -1579 -763 -1576 -747
rect -1568 -751 -1565 -739
rect -1521 -752 -1518 -737
rect -955 -752 -952 -736
rect -944 -740 -941 -728
rect -897 -741 -894 -726
rect -800 -732 -797 -728
rect -944 -752 -941 -744
rect -1568 -763 -1565 -755
rect -2474 -791 -2471 -788
rect -2463 -791 -2460 -788
rect -2261 -787 -2258 -772
rect -1734 -775 -1731 -772
rect -1723 -775 -1720 -772
rect -1521 -771 -1518 -756
rect -897 -760 -894 -745
rect -800 -752 -797 -736
rect -789 -740 -786 -728
rect -742 -741 -739 -726
rect -275 -727 -272 -723
rect -264 -727 -261 -723
rect -217 -727 -214 -724
rect -120 -727 -117 -723
rect -109 -727 -106 -723
rect -62 -727 -59 -724
rect -275 -738 -272 -734
rect -789 -752 -786 -744
rect -955 -764 -952 -761
rect -944 -764 -941 -761
rect -742 -760 -739 -745
rect -800 -764 -797 -761
rect -789 -764 -786 -761
rect -525 -761 -522 -757
rect -514 -761 -511 -757
rect -275 -758 -272 -742
rect -264 -746 -261 -734
rect -217 -747 -214 -732
rect -120 -738 -117 -734
rect -264 -758 -261 -750
rect -1579 -775 -1576 -772
rect -1568 -775 -1565 -772
rect -1304 -772 -1301 -768
rect -1293 -772 -1290 -768
rect -897 -769 -894 -765
rect -742 -769 -739 -765
rect -217 -766 -214 -751
rect -120 -758 -117 -742
rect -109 -746 -106 -734
rect -62 -747 -59 -732
rect -109 -758 -106 -750
rect -525 -772 -522 -768
rect -1676 -780 -1673 -776
rect -1521 -780 -1518 -776
rect -1304 -783 -1301 -779
rect -2319 -791 -2316 -788
rect -2308 -791 -2305 -788
rect -2044 -788 -2041 -784
rect -2033 -788 -2030 -784
rect -2416 -796 -2413 -792
rect -2261 -796 -2258 -792
rect -2044 -799 -2041 -795
rect -2044 -819 -2041 -803
rect -2033 -807 -2030 -795
rect -1304 -803 -1301 -787
rect -1293 -791 -1290 -779
rect -525 -792 -522 -776
rect -514 -780 -511 -768
rect -275 -770 -272 -767
rect -264 -770 -261 -767
rect -62 -766 -59 -751
rect -120 -770 -117 -767
rect -109 -770 -106 -767
rect 155 -767 158 -763
rect 166 -767 169 -763
rect -217 -775 -214 -771
rect -62 -775 -59 -771
rect 155 -778 158 -774
rect -514 -792 -511 -784
rect -1293 -803 -1290 -795
rect 155 -798 158 -782
rect 166 -786 169 -774
rect 166 -798 169 -790
rect -2033 -819 -2030 -811
rect -525 -804 -522 -801
rect -514 -804 -511 -801
rect 155 -810 158 -807
rect 166 -810 169 -807
rect -1304 -815 -1301 -812
rect -1293 -815 -1290 -812
rect -2044 -831 -2041 -828
rect -2033 -831 -2030 -828
<< ndiffusion >>
rect -2351 -525 -2348 -524
rect -2349 -529 -2348 -525
rect -2346 -525 -2342 -524
rect -2332 -525 -2329 -524
rect -2346 -529 -2344 -525
rect -2330 -529 -2329 -525
rect -2327 -525 -2321 -524
rect -2327 -529 -2325 -525
rect -2309 -525 -2304 -524
rect -2305 -529 -2304 -525
rect -2302 -525 -2299 -524
rect -2290 -525 -2285 -524
rect -2302 -529 -2300 -525
rect -2286 -529 -2285 -525
rect -2283 -525 -2279 -524
rect -2283 -529 -2281 -525
rect -1611 -509 -1608 -508
rect -1609 -513 -1608 -509
rect -1606 -509 -1602 -508
rect -1592 -509 -1589 -508
rect -1606 -513 -1604 -509
rect -1590 -513 -1589 -509
rect -1587 -509 -1581 -508
rect -1587 -513 -1585 -509
rect -1569 -509 -1564 -508
rect -1565 -513 -1564 -509
rect -1562 -509 -1559 -508
rect -1550 -509 -1545 -508
rect -1562 -513 -1560 -509
rect -1546 -513 -1545 -509
rect -1543 -509 -1539 -508
rect -1543 -513 -1541 -509
rect -832 -498 -829 -497
rect -830 -502 -829 -498
rect -827 -498 -823 -497
rect -813 -498 -810 -497
rect -827 -502 -825 -498
rect -811 -502 -810 -498
rect -808 -498 -802 -497
rect -808 -502 -806 -498
rect -790 -498 -785 -497
rect -786 -502 -785 -498
rect -783 -498 -780 -497
rect -771 -498 -766 -497
rect -783 -502 -781 -498
rect -767 -502 -766 -498
rect -764 -498 -760 -497
rect -764 -502 -762 -498
rect -152 -504 -149 -503
rect -150 -508 -149 -504
rect -147 -504 -143 -503
rect -133 -504 -130 -503
rect -147 -508 -145 -504
rect -131 -508 -130 -504
rect -128 -504 -122 -503
rect -128 -508 -126 -504
rect -110 -504 -105 -503
rect -106 -508 -105 -504
rect -103 -504 -100 -503
rect -91 -504 -86 -503
rect -103 -508 -101 -504
rect -87 -508 -86 -504
rect -84 -504 -80 -503
rect -84 -508 -82 -504
rect -2477 -691 -2474 -690
rect -2475 -695 -2474 -691
rect -2472 -691 -2468 -690
rect -2458 -691 -2455 -690
rect -2472 -695 -2470 -691
rect -2456 -695 -2455 -691
rect -2453 -691 -2447 -690
rect -2453 -695 -2451 -691
rect -2435 -691 -2430 -690
rect -2431 -695 -2430 -691
rect -2428 -691 -2425 -690
rect -2416 -691 -2411 -690
rect -2428 -695 -2426 -691
rect -2412 -695 -2411 -691
rect -2409 -691 -2405 -690
rect -2409 -695 -2407 -691
rect -2272 -687 -2269 -686
rect -2270 -691 -2269 -687
rect -2267 -687 -2263 -686
rect -2253 -687 -2250 -686
rect -2267 -691 -2265 -687
rect -2251 -691 -2250 -687
rect -2248 -687 -2242 -686
rect -2248 -691 -2246 -687
rect -2230 -687 -2225 -686
rect -2226 -691 -2225 -687
rect -2223 -687 -2220 -686
rect -2211 -687 -2206 -686
rect -2223 -691 -2221 -687
rect -2207 -691 -2206 -687
rect -2204 -687 -2200 -686
rect -2204 -691 -2202 -687
rect -1737 -675 -1734 -674
rect -1735 -679 -1734 -675
rect -1732 -675 -1728 -674
rect -1718 -675 -1715 -674
rect -1732 -679 -1730 -675
rect -1716 -679 -1715 -675
rect -1713 -675 -1707 -674
rect -1713 -679 -1711 -675
rect -1695 -675 -1690 -674
rect -1691 -679 -1690 -675
rect -1688 -675 -1685 -674
rect -1676 -675 -1671 -674
rect -1688 -679 -1686 -675
rect -1672 -679 -1671 -675
rect -1669 -675 -1665 -674
rect -1669 -679 -1667 -675
rect -1532 -671 -1529 -670
rect -1530 -675 -1529 -671
rect -1527 -671 -1523 -670
rect -1513 -671 -1510 -670
rect -1527 -675 -1525 -671
rect -1511 -675 -1510 -671
rect -1508 -671 -1502 -670
rect -1508 -675 -1506 -671
rect -1490 -671 -1485 -670
rect -1486 -675 -1485 -671
rect -1483 -671 -1480 -670
rect -1471 -671 -1466 -670
rect -1483 -675 -1481 -671
rect -1467 -675 -1466 -671
rect -1464 -671 -1460 -670
rect -1464 -675 -1462 -671
rect -2103 -728 -2101 -724
rect -2107 -733 -2101 -728
rect -2098 -733 -2090 -724
rect -2087 -728 -2084 -724
rect -2080 -728 -2079 -724
rect -958 -664 -955 -663
rect -956 -668 -955 -664
rect -953 -664 -949 -663
rect -939 -664 -936 -663
rect -953 -668 -951 -664
rect -937 -668 -936 -664
rect -934 -664 -928 -663
rect -934 -668 -932 -664
rect -916 -664 -911 -663
rect -912 -668 -911 -664
rect -909 -664 -906 -663
rect -897 -664 -892 -663
rect -909 -668 -907 -664
rect -893 -668 -892 -664
rect -890 -664 -886 -663
rect -890 -668 -888 -664
rect -753 -660 -750 -659
rect -751 -664 -750 -660
rect -748 -660 -744 -659
rect -734 -660 -731 -659
rect -748 -664 -746 -660
rect -732 -664 -731 -660
rect -729 -660 -723 -659
rect -729 -664 -727 -660
rect -711 -660 -706 -659
rect -707 -664 -706 -660
rect -704 -660 -701 -659
rect -692 -660 -687 -659
rect -704 -664 -702 -660
rect -688 -664 -687 -660
rect -685 -660 -681 -659
rect -685 -664 -683 -660
rect -1363 -712 -1361 -708
rect -1367 -717 -1361 -712
rect -1358 -717 -1350 -708
rect -1347 -712 -1344 -708
rect -1340 -712 -1339 -708
rect -584 -701 -582 -697
rect -588 -706 -582 -701
rect -579 -706 -571 -697
rect -568 -701 -565 -697
rect -561 -701 -560 -697
rect -278 -670 -275 -669
rect -276 -674 -275 -670
rect -273 -670 -269 -669
rect -259 -670 -256 -669
rect -273 -674 -271 -670
rect -257 -674 -256 -670
rect -254 -670 -248 -669
rect -254 -674 -252 -670
rect -236 -670 -231 -669
rect -232 -674 -231 -670
rect -229 -670 -226 -669
rect -217 -670 -212 -669
rect -229 -674 -227 -670
rect -213 -674 -212 -670
rect -210 -670 -206 -669
rect -210 -674 -208 -670
rect -73 -666 -70 -665
rect -71 -670 -70 -666
rect -68 -666 -64 -665
rect -54 -666 -51 -665
rect -68 -670 -66 -666
rect -52 -670 -51 -666
rect -49 -666 -43 -665
rect -49 -670 -47 -666
rect -31 -666 -26 -665
rect -27 -670 -26 -666
rect -24 -666 -21 -665
rect -12 -666 -7 -665
rect -24 -670 -22 -666
rect -8 -670 -7 -666
rect -5 -666 -1 -665
rect -5 -670 -3 -666
rect -568 -706 -560 -701
rect -506 -702 -504 -698
rect -510 -707 -504 -702
rect -501 -707 -493 -698
rect -490 -702 -487 -698
rect -483 -702 -482 -698
rect -490 -707 -482 -702
rect 96 -707 98 -703
rect -1347 -717 -1339 -712
rect -1285 -713 -1283 -709
rect -1289 -718 -1283 -713
rect -1280 -718 -1272 -709
rect -1269 -713 -1266 -709
rect -1262 -713 -1261 -709
rect -1269 -718 -1261 -713
rect 92 -712 98 -707
rect 101 -712 109 -703
rect 112 -707 115 -703
rect 119 -707 120 -703
rect 112 -712 120 -707
rect 174 -708 176 -704
rect 170 -713 176 -708
rect 179 -713 187 -704
rect 190 -708 193 -704
rect 197 -708 198 -704
rect 190 -713 198 -708
rect -2087 -733 -2079 -728
rect -2025 -729 -2023 -725
rect -2029 -734 -2023 -729
rect -2020 -734 -2012 -725
rect -2009 -729 -2006 -725
rect -2002 -729 -2001 -725
rect -2009 -734 -2001 -729
rect -2476 -783 -2474 -779
rect -2480 -788 -2474 -783
rect -2471 -788 -2463 -779
rect -2460 -783 -2457 -779
rect -2453 -783 -2452 -779
rect -2460 -788 -2452 -783
rect -1736 -767 -1734 -763
rect -1740 -772 -1734 -767
rect -1731 -772 -1723 -763
rect -1720 -767 -1717 -763
rect -1713 -767 -1712 -763
rect -1720 -772 -1712 -767
rect -1581 -767 -1579 -763
rect -2321 -783 -2319 -779
rect -2419 -792 -2416 -787
rect -2413 -792 -2409 -787
rect -2325 -788 -2319 -783
rect -2316 -788 -2308 -779
rect -2305 -783 -2302 -779
rect -2298 -783 -2297 -779
rect -2305 -788 -2297 -783
rect -1679 -776 -1676 -771
rect -1673 -776 -1669 -771
rect -1585 -772 -1579 -767
rect -1576 -772 -1568 -763
rect -1565 -767 -1562 -763
rect -1558 -767 -1557 -763
rect -1565 -772 -1557 -767
rect -957 -756 -955 -752
rect -961 -761 -955 -756
rect -952 -761 -944 -752
rect -941 -756 -938 -752
rect -934 -756 -933 -752
rect -941 -761 -933 -756
rect -802 -756 -800 -752
rect -900 -765 -897 -760
rect -894 -765 -890 -760
rect -806 -761 -800 -756
rect -797 -761 -789 -752
rect -786 -756 -783 -752
rect -779 -756 -778 -752
rect -786 -761 -778 -756
rect -745 -765 -742 -760
rect -739 -765 -735 -760
rect -1524 -776 -1521 -771
rect -1518 -776 -1514 -771
rect -277 -762 -275 -758
rect -281 -767 -275 -762
rect -272 -767 -264 -758
rect -261 -762 -258 -758
rect -254 -762 -253 -758
rect -261 -767 -253 -762
rect -122 -762 -120 -758
rect -2264 -792 -2261 -787
rect -2258 -792 -2254 -787
rect -220 -771 -217 -766
rect -214 -771 -210 -766
rect -126 -767 -120 -762
rect -117 -767 -109 -758
rect -106 -762 -103 -758
rect -99 -762 -98 -758
rect -106 -767 -98 -762
rect -65 -771 -62 -766
rect -59 -771 -55 -766
rect -527 -796 -525 -792
rect -531 -801 -525 -796
rect -522 -801 -514 -792
rect -511 -796 -508 -792
rect -504 -796 -503 -792
rect -511 -801 -503 -796
rect -1306 -807 -1304 -803
rect -1310 -812 -1304 -807
rect -1301 -812 -1293 -803
rect -1290 -807 -1287 -803
rect -1283 -807 -1282 -803
rect 153 -802 155 -798
rect 149 -807 155 -802
rect 158 -807 166 -798
rect 169 -802 172 -798
rect 176 -802 177 -798
rect 169 -807 177 -802
rect -1290 -812 -1282 -807
rect -2046 -823 -2044 -819
rect -2050 -828 -2044 -823
rect -2041 -828 -2033 -819
rect -2030 -823 -2027 -819
rect -2023 -823 -2022 -819
rect -2030 -828 -2022 -823
<< pdiffusion >>
rect -2353 -494 -2348 -493
rect -2349 -498 -2348 -494
rect -2346 -494 -2340 -493
rect -2346 -498 -2344 -494
rect -2334 -494 -2329 -493
rect -2330 -498 -2329 -494
rect -2327 -494 -2321 -493
rect -2327 -498 -2325 -494
rect -2309 -494 -2304 -493
rect -2305 -498 -2304 -494
rect -2302 -494 -2296 -493
rect -2302 -498 -2300 -494
rect -2290 -494 -2285 -493
rect -2286 -498 -2285 -494
rect -2283 -494 -2277 -493
rect -2283 -498 -2281 -494
rect -1613 -478 -1608 -477
rect -1609 -482 -1608 -478
rect -1606 -478 -1600 -477
rect -1606 -482 -1604 -478
rect -1594 -478 -1589 -477
rect -1590 -482 -1589 -478
rect -1587 -478 -1581 -477
rect -1587 -482 -1585 -478
rect -1569 -478 -1564 -477
rect -1565 -482 -1564 -478
rect -1562 -478 -1556 -477
rect -1562 -482 -1560 -478
rect -1550 -478 -1545 -477
rect -1546 -482 -1545 -478
rect -1543 -478 -1537 -477
rect -1543 -482 -1541 -478
rect -834 -467 -829 -466
rect -830 -471 -829 -467
rect -827 -467 -821 -466
rect -827 -471 -825 -467
rect -815 -467 -810 -466
rect -811 -471 -810 -467
rect -808 -467 -802 -466
rect -808 -471 -806 -467
rect -790 -467 -785 -466
rect -786 -471 -785 -467
rect -783 -467 -777 -466
rect -783 -471 -781 -467
rect -771 -467 -766 -466
rect -767 -471 -766 -467
rect -764 -467 -758 -466
rect -764 -471 -762 -467
rect -154 -473 -149 -472
rect -150 -477 -149 -473
rect -147 -473 -141 -472
rect -147 -477 -145 -473
rect -135 -473 -130 -472
rect -131 -477 -130 -473
rect -128 -473 -122 -472
rect -128 -477 -126 -473
rect -110 -473 -105 -472
rect -106 -477 -105 -473
rect -103 -473 -97 -472
rect -103 -477 -101 -473
rect -91 -473 -86 -472
rect -87 -477 -86 -473
rect -84 -473 -78 -472
rect -84 -477 -82 -473
rect -2479 -660 -2474 -659
rect -2475 -664 -2474 -660
rect -2472 -660 -2466 -659
rect -2472 -664 -2470 -660
rect -2460 -660 -2455 -659
rect -2456 -664 -2455 -660
rect -2453 -660 -2447 -659
rect -2453 -664 -2451 -660
rect -2435 -660 -2430 -659
rect -2431 -664 -2430 -660
rect -2428 -660 -2422 -659
rect -2428 -664 -2426 -660
rect -2416 -660 -2411 -659
rect -2412 -664 -2411 -660
rect -2409 -660 -2403 -659
rect -2409 -664 -2407 -660
rect -2274 -656 -2269 -655
rect -2270 -660 -2269 -656
rect -2267 -656 -2261 -655
rect -2267 -660 -2265 -656
rect -2255 -656 -2250 -655
rect -2251 -660 -2250 -656
rect -2248 -656 -2242 -655
rect -2248 -660 -2246 -656
rect -2230 -656 -2225 -655
rect -2226 -660 -2225 -656
rect -2223 -656 -2217 -655
rect -2223 -660 -2221 -656
rect -2211 -656 -2206 -655
rect -2207 -660 -2206 -656
rect -2204 -656 -2198 -655
rect -2204 -660 -2202 -656
rect -2104 -697 -2101 -693
rect -2108 -700 -2101 -697
rect -2098 -697 -2095 -693
rect -2091 -697 -2090 -693
rect -2098 -700 -2090 -697
rect -2087 -697 -2084 -693
rect -1739 -644 -1734 -643
rect -1735 -648 -1734 -644
rect -1732 -644 -1726 -643
rect -1732 -648 -1730 -644
rect -1720 -644 -1715 -643
rect -1716 -648 -1715 -644
rect -1713 -644 -1707 -643
rect -1713 -648 -1711 -644
rect -1695 -644 -1690 -643
rect -1691 -648 -1690 -644
rect -1688 -644 -1682 -643
rect -1688 -648 -1686 -644
rect -1676 -644 -1671 -643
rect -1672 -648 -1671 -644
rect -1669 -644 -1663 -643
rect -1669 -648 -1667 -644
rect -1534 -640 -1529 -639
rect -1530 -644 -1529 -640
rect -1527 -640 -1521 -639
rect -1527 -644 -1525 -640
rect -1515 -640 -1510 -639
rect -1511 -644 -1510 -640
rect -1508 -640 -1502 -639
rect -1508 -644 -1506 -640
rect -1490 -640 -1485 -639
rect -1486 -644 -1485 -640
rect -1483 -640 -1477 -639
rect -1483 -644 -1481 -640
rect -1471 -640 -1466 -639
rect -1467 -644 -1466 -640
rect -1464 -640 -1458 -639
rect -1464 -644 -1462 -640
rect -1364 -681 -1361 -677
rect -1368 -684 -1361 -681
rect -1358 -681 -1355 -677
rect -1351 -681 -1350 -677
rect -1358 -684 -1350 -681
rect -1347 -681 -1344 -677
rect -1347 -684 -1340 -681
rect -1286 -682 -1283 -678
rect -2087 -700 -2080 -697
rect -2026 -698 -2023 -694
rect -2030 -701 -2023 -698
rect -2020 -698 -2017 -694
rect -2013 -698 -2012 -694
rect -2020 -701 -2012 -698
rect -2009 -698 -2006 -694
rect -2009 -701 -2002 -698
rect -1290 -685 -1283 -682
rect -1280 -682 -1277 -678
rect -1273 -682 -1272 -678
rect -1280 -685 -1272 -682
rect -1269 -682 -1266 -678
rect -960 -633 -955 -632
rect -956 -637 -955 -633
rect -953 -633 -947 -632
rect -953 -637 -951 -633
rect -941 -633 -936 -632
rect -937 -637 -936 -633
rect -934 -633 -928 -632
rect -934 -637 -932 -633
rect -916 -633 -911 -632
rect -912 -637 -911 -633
rect -909 -633 -903 -632
rect -909 -637 -907 -633
rect -897 -633 -892 -632
rect -893 -637 -892 -633
rect -890 -633 -884 -632
rect -890 -637 -888 -633
rect -755 -629 -750 -628
rect -751 -633 -750 -629
rect -748 -629 -742 -628
rect -748 -633 -746 -629
rect -736 -629 -731 -628
rect -732 -633 -731 -629
rect -729 -629 -723 -628
rect -729 -633 -727 -629
rect -711 -629 -706 -628
rect -707 -633 -706 -629
rect -704 -629 -698 -628
rect -704 -633 -702 -629
rect -692 -629 -687 -628
rect -688 -633 -687 -629
rect -685 -629 -679 -628
rect -685 -633 -683 -629
rect -585 -670 -582 -666
rect -589 -673 -582 -670
rect -579 -670 -576 -666
rect -572 -670 -571 -666
rect -579 -673 -571 -670
rect -568 -670 -565 -666
rect -568 -673 -561 -670
rect -507 -671 -504 -667
rect -1269 -685 -1262 -682
rect -511 -674 -504 -671
rect -501 -671 -498 -667
rect -494 -671 -493 -667
rect -501 -674 -493 -671
rect -490 -671 -487 -667
rect -490 -674 -483 -671
rect -280 -639 -275 -638
rect -276 -643 -275 -639
rect -273 -639 -267 -638
rect -273 -643 -271 -639
rect -261 -639 -256 -638
rect -257 -643 -256 -639
rect -254 -639 -248 -638
rect -254 -643 -252 -639
rect -236 -639 -231 -638
rect -232 -643 -231 -639
rect -229 -639 -223 -638
rect -229 -643 -227 -639
rect -217 -639 -212 -638
rect -213 -643 -212 -639
rect -210 -639 -204 -638
rect -210 -643 -208 -639
rect -75 -635 -70 -634
rect -71 -639 -70 -635
rect -68 -635 -62 -634
rect -68 -639 -66 -635
rect -56 -635 -51 -634
rect -52 -639 -51 -635
rect -49 -635 -43 -634
rect -49 -639 -47 -635
rect -31 -635 -26 -634
rect -27 -639 -26 -635
rect -24 -635 -18 -634
rect -24 -639 -22 -635
rect -12 -635 -7 -634
rect -8 -639 -7 -635
rect -5 -635 1 -634
rect -5 -639 -3 -635
rect 95 -676 98 -672
rect 91 -679 98 -676
rect 101 -676 104 -672
rect 108 -676 109 -672
rect 101 -679 109 -676
rect 112 -676 115 -672
rect 112 -679 119 -676
rect 173 -677 176 -673
rect 169 -680 176 -677
rect 179 -677 182 -673
rect 186 -677 187 -673
rect 179 -680 187 -677
rect 190 -677 193 -673
rect 190 -680 197 -677
rect -958 -725 -955 -721
rect -962 -728 -955 -725
rect -952 -725 -949 -721
rect -945 -725 -944 -721
rect -952 -728 -944 -725
rect -941 -725 -938 -721
rect -941 -728 -934 -725
rect -901 -726 -897 -721
rect -894 -726 -890 -721
rect -886 -726 -884 -721
rect -803 -725 -800 -721
rect -1737 -736 -1734 -732
rect -1741 -739 -1734 -736
rect -1731 -736 -1728 -732
rect -1724 -736 -1723 -732
rect -1731 -739 -1723 -736
rect -1720 -736 -1717 -732
rect -1720 -739 -1713 -736
rect -1680 -737 -1676 -732
rect -1673 -737 -1669 -732
rect -1665 -737 -1663 -732
rect -1582 -736 -1579 -732
rect -2477 -752 -2474 -748
rect -2481 -755 -2474 -752
rect -2471 -752 -2468 -748
rect -2464 -752 -2463 -748
rect -2471 -755 -2463 -752
rect -2460 -752 -2457 -748
rect -2460 -755 -2453 -752
rect -2420 -753 -2416 -748
rect -2413 -753 -2409 -748
rect -2405 -753 -2403 -748
rect -2322 -752 -2319 -748
rect -2326 -755 -2319 -752
rect -2316 -752 -2313 -748
rect -2309 -752 -2308 -748
rect -2316 -755 -2308 -752
rect -2305 -752 -2302 -748
rect -2305 -755 -2298 -752
rect -2265 -753 -2261 -748
rect -2258 -753 -2254 -748
rect -2250 -753 -2248 -748
rect -1586 -739 -1579 -736
rect -1576 -736 -1573 -732
rect -1569 -736 -1568 -732
rect -1576 -739 -1568 -736
rect -1565 -736 -1562 -732
rect -1565 -739 -1558 -736
rect -1525 -737 -1521 -732
rect -1518 -737 -1514 -732
rect -1510 -737 -1508 -732
rect -807 -728 -800 -725
rect -797 -725 -794 -721
rect -790 -725 -789 -721
rect -797 -728 -789 -725
rect -786 -725 -783 -721
rect -786 -728 -779 -725
rect -746 -726 -742 -721
rect -739 -726 -735 -721
rect -731 -726 -729 -721
rect -278 -731 -275 -727
rect -282 -734 -275 -731
rect -272 -731 -269 -727
rect -265 -731 -264 -727
rect -272 -734 -264 -731
rect -261 -731 -258 -727
rect -261 -734 -254 -731
rect -221 -732 -217 -727
rect -214 -732 -210 -727
rect -206 -732 -204 -727
rect -123 -731 -120 -727
rect -127 -734 -120 -731
rect -117 -731 -114 -727
rect -110 -731 -109 -727
rect -117 -734 -109 -731
rect -106 -731 -103 -727
rect -106 -734 -99 -731
rect -66 -732 -62 -727
rect -59 -732 -55 -727
rect -51 -732 -49 -727
rect -528 -765 -525 -761
rect -532 -768 -525 -765
rect -522 -765 -519 -761
rect -515 -765 -514 -761
rect -522 -768 -514 -765
rect -511 -765 -508 -761
rect -511 -768 -504 -765
rect -1307 -776 -1304 -772
rect -1311 -779 -1304 -776
rect -1301 -776 -1298 -772
rect -1294 -776 -1293 -772
rect -1301 -779 -1293 -776
rect -1290 -776 -1287 -772
rect -1290 -779 -1283 -776
rect -2047 -792 -2044 -788
rect -2051 -795 -2044 -792
rect -2041 -792 -2038 -788
rect -2034 -792 -2033 -788
rect -2041 -795 -2033 -792
rect -2030 -792 -2027 -788
rect -2030 -795 -2023 -792
rect 152 -771 155 -767
rect 148 -774 155 -771
rect 158 -771 161 -767
rect 165 -771 166 -767
rect 158 -774 166 -771
rect 169 -771 172 -767
rect 169 -774 176 -771
<< metal1 >>
rect -1232 -369 -1079 -365
rect -1972 -385 -1897 -381
rect -2353 -470 -2312 -466
rect -2353 -494 -2349 -470
rect -2353 -525 -2349 -498
rect -2344 -494 -2340 -473
rect -2336 -477 -2320 -473
rect -2325 -494 -2321 -477
rect -2344 -525 -2340 -498
rect -2334 -525 -2330 -498
rect -2325 -525 -2321 -498
rect -2317 -510 -2313 -470
rect -2309 -481 -2285 -478
rect -2309 -482 -2286 -481
rect -2309 -494 -2305 -482
rect -2290 -494 -2286 -482
rect -2317 -514 -2307 -510
rect -2300 -518 -2296 -498
rect -2281 -510 -2277 -498
rect -2290 -514 -2288 -510
rect -2281 -514 -2278 -510
rect -2317 -522 -2296 -518
rect -2334 -532 -2330 -529
rect -2317 -532 -2313 -522
rect -2300 -525 -2296 -522
rect -2281 -525 -2277 -514
rect -2334 -536 -2313 -532
rect -2309 -532 -2305 -529
rect -2290 -531 -2286 -529
rect -2291 -532 -2286 -531
rect -2309 -536 -2286 -532
rect -2448 -632 -2444 -630
rect -2274 -632 -2244 -628
rect -2240 -632 -2234 -628
rect -2479 -636 -2439 -632
rect -2479 -660 -2475 -636
rect -2479 -691 -2475 -664
rect -2470 -643 -2451 -639
rect -2470 -644 -2465 -643
rect -2470 -660 -2466 -644
rect -2451 -660 -2447 -643
rect -2470 -691 -2466 -664
rect -2460 -691 -2456 -664
rect -2451 -691 -2447 -664
rect -2443 -675 -2439 -636
rect -2435 -648 -2412 -644
rect -2435 -660 -2431 -648
rect -2416 -660 -2412 -648
rect -2274 -656 -2270 -632
rect -2443 -676 -2438 -675
rect -2443 -680 -2433 -676
rect -2426 -684 -2422 -664
rect -2407 -676 -2403 -664
rect -2417 -683 -2414 -677
rect -2407 -680 -2404 -676
rect -2443 -688 -2422 -684
rect -2460 -698 -2456 -695
rect -2443 -698 -2439 -688
rect -2426 -691 -2422 -688
rect -2407 -691 -2403 -680
rect -2274 -687 -2270 -660
rect -2265 -639 -2242 -635
rect -2265 -656 -2261 -639
rect -2246 -656 -2242 -639
rect -2265 -687 -2261 -660
rect -2255 -687 -2251 -660
rect -2246 -687 -2242 -660
rect -2238 -672 -2234 -632
rect -2221 -639 -2217 -638
rect -2221 -640 -2214 -639
rect -2230 -644 -2207 -640
rect -2230 -656 -2226 -644
rect -2211 -656 -2207 -644
rect -2238 -676 -2228 -672
rect -2221 -680 -2217 -660
rect -2202 -672 -2198 -660
rect -2213 -679 -2209 -672
rect -2202 -676 -2199 -672
rect -2238 -684 -2217 -680
rect -2210 -683 -2209 -679
rect -2460 -702 -2439 -698
rect -2255 -694 -2251 -691
rect -2238 -694 -2234 -684
rect -2221 -687 -2217 -684
rect -2202 -687 -2198 -676
rect -2098 -683 -2086 -682
rect -2435 -698 -2431 -695
rect -2418 -697 -2412 -695
rect -2419 -698 -2412 -697
rect -2255 -698 -2234 -694
rect -2108 -684 -2015 -683
rect -2108 -687 -2002 -684
rect -2230 -694 -2226 -691
rect -2211 -692 -2207 -691
rect -2214 -694 -2207 -692
rect -2230 -695 -2207 -694
rect -2231 -698 -2207 -695
rect -2108 -693 -2104 -687
rect -2084 -693 -2080 -687
rect -2030 -688 -2002 -687
rect -2030 -694 -2026 -688
rect -2006 -694 -2002 -688
rect -2435 -702 -2412 -698
rect -2095 -704 -2091 -697
rect -2134 -708 -2102 -704
rect -2095 -707 -2080 -704
rect -2017 -705 -2013 -698
rect -2316 -738 -2304 -737
rect -2481 -742 -2421 -738
rect -2417 -742 -2392 -738
rect -2326 -742 -2266 -738
rect -2262 -742 -2237 -738
rect -2481 -748 -2477 -742
rect -2457 -748 -2453 -742
rect -2424 -748 -2421 -742
rect -2326 -748 -2322 -742
rect -2302 -748 -2298 -742
rect -2468 -759 -2464 -752
rect -2269 -748 -2266 -742
rect -2486 -763 -2475 -759
rect -2468 -762 -2453 -759
rect -2457 -765 -2453 -762
rect -2482 -771 -2464 -767
rect -2457 -768 -2452 -765
rect -2408 -768 -2405 -753
rect -2313 -759 -2309 -752
rect -2327 -763 -2320 -759
rect -2313 -762 -2298 -759
rect -2302 -765 -2298 -762
rect -2457 -772 -2417 -768
rect -2408 -771 -2382 -768
rect -2328 -771 -2309 -767
rect -2302 -768 -2297 -765
rect -2253 -767 -2250 -753
rect -2457 -779 -2453 -772
rect -2480 -792 -2476 -783
rect -2408 -787 -2405 -771
rect -2480 -793 -2448 -792
rect -2424 -793 -2420 -792
rect -2480 -795 -2420 -793
rect -2452 -796 -2420 -795
rect -2385 -819 -2382 -771
rect -2302 -772 -2262 -768
rect -2253 -771 -2248 -767
rect -2302 -779 -2298 -772
rect -2325 -792 -2321 -783
rect -2253 -787 -2250 -771
rect -2325 -795 -2279 -792
rect -2298 -796 -2278 -795
rect -2269 -796 -2265 -792
rect -2298 -797 -2265 -796
rect -2297 -799 -2265 -797
rect -2134 -819 -2131 -708
rect -2109 -712 -2106 -708
rect -2084 -710 -2080 -707
rect -2032 -709 -2024 -705
rect -2017 -708 -2002 -705
rect -2109 -716 -2091 -712
rect -2084 -713 -2079 -710
rect -2032 -713 -2028 -709
rect -2006 -711 -2002 -708
rect -2006 -713 -2001 -711
rect -2084 -717 -2072 -713
rect -2032 -717 -2013 -713
rect -2006 -716 -1994 -713
rect -2084 -724 -2080 -717
rect -2107 -737 -2103 -728
rect -2107 -740 -2078 -737
rect -2100 -742 -2090 -740
rect -2075 -807 -2072 -717
rect -2006 -725 -2002 -716
rect -2029 -738 -2025 -729
rect -2029 -741 -2000 -738
rect -2020 -743 -2012 -741
rect -1997 -767 -1994 -716
rect -2069 -770 -1994 -767
rect -2069 -799 -2065 -770
rect -2044 -778 -2033 -775
rect -2051 -782 -2023 -778
rect -2051 -788 -2047 -782
rect -2027 -788 -2023 -782
rect -2038 -799 -2034 -792
rect -2069 -803 -2045 -799
rect -2038 -802 -2023 -799
rect -2027 -805 -2023 -802
rect -2075 -811 -2034 -807
rect -2027 -808 -2010 -805
rect -2027 -809 -2015 -808
rect -2027 -819 -2023 -809
rect -2385 -822 -2131 -819
rect -2050 -832 -2046 -823
rect -2050 -835 -2021 -832
rect -2039 -837 -2028 -835
rect -1902 -878 -1898 -385
rect -1613 -454 -1572 -450
rect -1613 -478 -1609 -454
rect -1613 -509 -1609 -482
rect -1604 -478 -1600 -457
rect -1596 -461 -1580 -457
rect -1585 -478 -1581 -461
rect -1604 -509 -1600 -482
rect -1594 -509 -1590 -482
rect -1585 -509 -1581 -482
rect -1577 -494 -1573 -454
rect -1569 -465 -1545 -462
rect -1569 -466 -1546 -465
rect -1569 -478 -1565 -466
rect -1550 -478 -1546 -466
rect -1577 -498 -1567 -494
rect -1560 -502 -1556 -482
rect -1541 -494 -1537 -482
rect -1550 -498 -1548 -494
rect -1541 -498 -1538 -494
rect -1577 -506 -1556 -502
rect -1594 -516 -1590 -513
rect -1577 -516 -1573 -506
rect -1560 -509 -1556 -506
rect -1541 -509 -1537 -498
rect -1594 -520 -1573 -516
rect -1569 -516 -1565 -513
rect -1550 -515 -1546 -513
rect -1551 -516 -1546 -515
rect -1569 -520 -1546 -516
rect -1708 -616 -1704 -614
rect -1534 -616 -1504 -612
rect -1500 -616 -1494 -612
rect -1739 -620 -1699 -616
rect -1739 -644 -1735 -620
rect -1739 -675 -1735 -648
rect -1730 -627 -1711 -623
rect -1730 -628 -1725 -627
rect -1730 -644 -1726 -628
rect -1711 -644 -1707 -627
rect -1730 -675 -1726 -648
rect -1720 -675 -1716 -648
rect -1711 -675 -1707 -648
rect -1703 -659 -1699 -620
rect -1695 -632 -1672 -628
rect -1695 -644 -1691 -632
rect -1676 -644 -1672 -632
rect -1534 -640 -1530 -616
rect -1703 -660 -1698 -659
rect -1703 -664 -1693 -660
rect -1686 -668 -1682 -648
rect -1667 -660 -1663 -648
rect -1677 -667 -1674 -661
rect -1667 -664 -1664 -660
rect -1703 -672 -1682 -668
rect -1720 -682 -1716 -679
rect -1703 -682 -1699 -672
rect -1686 -675 -1682 -672
rect -1667 -675 -1663 -664
rect -1534 -671 -1530 -644
rect -1525 -623 -1502 -619
rect -1525 -640 -1521 -623
rect -1506 -640 -1502 -623
rect -1525 -671 -1521 -644
rect -1515 -671 -1511 -644
rect -1506 -671 -1502 -644
rect -1498 -656 -1494 -616
rect -1481 -623 -1477 -622
rect -1481 -624 -1474 -623
rect -1490 -628 -1467 -624
rect -1490 -640 -1486 -628
rect -1471 -640 -1467 -628
rect -1498 -660 -1488 -656
rect -1481 -664 -1477 -644
rect -1462 -656 -1458 -644
rect -1473 -663 -1469 -656
rect -1462 -660 -1459 -656
rect -1498 -668 -1477 -664
rect -1470 -667 -1469 -663
rect -1720 -686 -1699 -682
rect -1515 -678 -1511 -675
rect -1498 -678 -1494 -668
rect -1481 -671 -1477 -668
rect -1462 -671 -1458 -660
rect -1358 -667 -1346 -666
rect -1695 -682 -1691 -679
rect -1678 -681 -1672 -679
rect -1679 -682 -1672 -681
rect -1515 -682 -1494 -678
rect -1368 -668 -1275 -667
rect -1368 -671 -1262 -668
rect -1490 -678 -1486 -675
rect -1471 -676 -1467 -675
rect -1474 -678 -1467 -676
rect -1490 -679 -1467 -678
rect -1491 -682 -1467 -679
rect -1368 -677 -1364 -671
rect -1344 -677 -1340 -671
rect -1290 -672 -1262 -671
rect -1290 -678 -1286 -672
rect -1266 -678 -1262 -672
rect -1695 -686 -1672 -682
rect -1355 -688 -1351 -681
rect -1394 -692 -1362 -688
rect -1355 -691 -1340 -688
rect -1277 -689 -1273 -682
rect -1576 -722 -1564 -721
rect -1741 -726 -1681 -722
rect -1677 -726 -1652 -722
rect -1586 -726 -1526 -722
rect -1522 -726 -1497 -722
rect -1741 -732 -1737 -726
rect -1717 -732 -1713 -726
rect -1684 -732 -1681 -726
rect -1586 -732 -1582 -726
rect -1562 -732 -1558 -726
rect -1728 -743 -1724 -736
rect -1529 -732 -1526 -726
rect -1746 -747 -1735 -743
rect -1728 -746 -1713 -743
rect -1717 -749 -1713 -746
rect -1742 -755 -1724 -751
rect -1717 -752 -1712 -749
rect -1668 -752 -1665 -737
rect -1573 -743 -1569 -736
rect -1587 -747 -1580 -743
rect -1573 -746 -1558 -743
rect -1562 -749 -1558 -746
rect -1717 -756 -1677 -752
rect -1668 -755 -1642 -752
rect -1588 -755 -1569 -751
rect -1562 -752 -1557 -749
rect -1513 -751 -1510 -737
rect -1717 -763 -1713 -756
rect -1740 -776 -1736 -767
rect -1668 -771 -1665 -755
rect -1740 -777 -1708 -776
rect -1684 -777 -1680 -776
rect -1740 -779 -1680 -777
rect -1712 -780 -1680 -779
rect -1645 -803 -1642 -755
rect -1562 -756 -1522 -752
rect -1513 -755 -1508 -751
rect -1562 -763 -1558 -756
rect -1585 -776 -1581 -767
rect -1513 -771 -1510 -755
rect -1585 -779 -1539 -776
rect -1558 -780 -1538 -779
rect -1529 -780 -1525 -776
rect -1558 -781 -1525 -780
rect -1557 -783 -1525 -781
rect -1557 -784 -1497 -783
rect -1539 -789 -1497 -784
rect -1394 -803 -1391 -692
rect -1369 -696 -1366 -692
rect -1344 -694 -1340 -691
rect -1292 -693 -1284 -689
rect -1277 -692 -1262 -689
rect -1369 -700 -1351 -696
rect -1344 -697 -1339 -694
rect -1292 -697 -1288 -693
rect -1266 -695 -1262 -692
rect -1266 -697 -1261 -695
rect -1344 -701 -1332 -697
rect -1292 -701 -1273 -697
rect -1266 -700 -1254 -697
rect -1344 -708 -1340 -701
rect -1367 -721 -1363 -712
rect -1367 -724 -1338 -721
rect -1360 -726 -1350 -724
rect -1335 -791 -1332 -701
rect -1266 -709 -1262 -700
rect -1289 -722 -1285 -713
rect -1289 -725 -1260 -722
rect -1280 -727 -1272 -725
rect -1257 -751 -1254 -700
rect -1329 -754 -1254 -751
rect -1329 -783 -1325 -754
rect -1304 -762 -1293 -759
rect -1311 -766 -1283 -762
rect -1311 -772 -1307 -766
rect -1287 -772 -1283 -766
rect -1298 -783 -1294 -776
rect -1329 -787 -1305 -783
rect -1298 -786 -1283 -783
rect -1287 -789 -1283 -786
rect -1335 -795 -1294 -791
rect -1287 -793 -1262 -789
rect -1287 -803 -1283 -793
rect -1645 -806 -1391 -803
rect -1310 -816 -1306 -807
rect -1310 -819 -1281 -816
rect -1299 -821 -1288 -819
rect -1266 -878 -1262 -793
rect -1083 -851 -1079 -369
rect -834 -443 -793 -439
rect -834 -467 -830 -443
rect -834 -498 -830 -471
rect -825 -467 -821 -446
rect -817 -450 -801 -446
rect -806 -467 -802 -450
rect -825 -498 -821 -471
rect -815 -498 -811 -471
rect -806 -498 -802 -471
rect -798 -483 -794 -443
rect -154 -449 -113 -445
rect -790 -454 -766 -451
rect -790 -455 -767 -454
rect -790 -467 -786 -455
rect -771 -467 -767 -455
rect -798 -487 -788 -483
rect -781 -491 -777 -471
rect -762 -483 -758 -471
rect -154 -473 -150 -449
rect -771 -487 -769 -483
rect -762 -487 -759 -483
rect -798 -495 -777 -491
rect -815 -505 -811 -502
rect -798 -505 -794 -495
rect -781 -498 -777 -495
rect -762 -498 -758 -487
rect -815 -509 -794 -505
rect -790 -505 -786 -502
rect -771 -504 -767 -502
rect -772 -505 -767 -504
rect -790 -509 -767 -505
rect -154 -504 -150 -477
rect -145 -473 -141 -452
rect -137 -456 -121 -452
rect -126 -473 -122 -456
rect -145 -504 -141 -477
rect -135 -504 -131 -477
rect -126 -504 -122 -477
rect -118 -489 -114 -449
rect -110 -460 -86 -457
rect -110 -461 -87 -460
rect -110 -473 -106 -461
rect -91 -473 -87 -461
rect -118 -493 -108 -489
rect -101 -497 -97 -477
rect -82 -489 -78 -477
rect -91 -493 -89 -489
rect -82 -493 -79 -489
rect -118 -501 -97 -497
rect -135 -511 -131 -508
rect -118 -511 -114 -501
rect -101 -504 -97 -501
rect -82 -504 -78 -493
rect -135 -515 -114 -511
rect -110 -511 -106 -508
rect -91 -510 -87 -508
rect -92 -511 -87 -510
rect -110 -515 -87 -511
rect -929 -605 -925 -603
rect -755 -605 -725 -601
rect -721 -605 -715 -601
rect -960 -609 -920 -605
rect -960 -633 -956 -609
rect -960 -664 -956 -637
rect -951 -616 -932 -612
rect -951 -617 -946 -616
rect -951 -633 -947 -617
rect -932 -633 -928 -616
rect -951 -664 -947 -637
rect -941 -664 -937 -637
rect -932 -664 -928 -637
rect -924 -648 -920 -609
rect -916 -621 -893 -617
rect -916 -633 -912 -621
rect -897 -633 -893 -621
rect -755 -629 -751 -605
rect -924 -649 -919 -648
rect -924 -653 -914 -649
rect -907 -657 -903 -637
rect -888 -649 -884 -637
rect -898 -656 -895 -650
rect -888 -653 -885 -649
rect -924 -661 -903 -657
rect -941 -671 -937 -668
rect -924 -671 -920 -661
rect -907 -664 -903 -661
rect -888 -664 -884 -653
rect -755 -660 -751 -633
rect -746 -612 -723 -608
rect -746 -629 -742 -612
rect -727 -629 -723 -612
rect -746 -660 -742 -633
rect -736 -660 -732 -633
rect -727 -660 -723 -633
rect -719 -645 -715 -605
rect -249 -611 -245 -609
rect -75 -611 -45 -607
rect -41 -611 -35 -607
rect -702 -612 -698 -611
rect -702 -613 -695 -612
rect -711 -617 -688 -613
rect -711 -629 -707 -617
rect -692 -629 -688 -617
rect -280 -615 -240 -611
rect -719 -649 -709 -645
rect -702 -653 -698 -633
rect -683 -645 -679 -633
rect -280 -639 -276 -615
rect -694 -652 -690 -645
rect -683 -649 -680 -645
rect -719 -657 -698 -653
rect -691 -656 -690 -652
rect -941 -675 -920 -671
rect -736 -667 -732 -664
rect -719 -667 -715 -657
rect -702 -660 -698 -657
rect -683 -660 -679 -649
rect -579 -656 -567 -655
rect -916 -671 -912 -668
rect -899 -670 -893 -668
rect -900 -671 -893 -670
rect -736 -671 -715 -667
rect -589 -657 -496 -656
rect -589 -660 -483 -657
rect -711 -667 -707 -664
rect -692 -665 -688 -664
rect -695 -667 -688 -665
rect -711 -668 -688 -667
rect -712 -671 -688 -668
rect -589 -666 -585 -660
rect -565 -666 -561 -660
rect -511 -661 -483 -660
rect -511 -667 -507 -661
rect -487 -667 -483 -661
rect -916 -675 -893 -671
rect -576 -677 -572 -670
rect -280 -670 -276 -643
rect -615 -681 -583 -677
rect -576 -680 -561 -677
rect -498 -678 -494 -671
rect -271 -622 -252 -618
rect -271 -623 -266 -622
rect -271 -639 -267 -623
rect -252 -639 -248 -622
rect -271 -670 -267 -643
rect -261 -670 -257 -643
rect -252 -670 -248 -643
rect -244 -654 -240 -615
rect -236 -627 -213 -623
rect -236 -639 -232 -627
rect -217 -639 -213 -627
rect -75 -635 -71 -611
rect -244 -655 -239 -654
rect -244 -659 -234 -655
rect -227 -663 -223 -643
rect -208 -655 -204 -643
rect -218 -662 -215 -656
rect -208 -659 -205 -655
rect -244 -667 -223 -663
rect -261 -677 -257 -674
rect -244 -677 -240 -667
rect -227 -670 -223 -667
rect -208 -670 -204 -659
rect -75 -666 -71 -639
rect -66 -618 -43 -614
rect -66 -635 -62 -618
rect -47 -635 -43 -618
rect -66 -666 -62 -639
rect -56 -666 -52 -639
rect -47 -666 -43 -639
rect -39 -651 -35 -611
rect -22 -618 -18 -617
rect -22 -619 -15 -618
rect -31 -623 -8 -619
rect -31 -635 -27 -623
rect -12 -635 -8 -623
rect -39 -655 -29 -651
rect -22 -659 -18 -639
rect -3 -651 1 -639
rect -13 -655 -10 -651
rect -3 -655 0 -651
rect -39 -663 -18 -659
rect -797 -711 -785 -710
rect -962 -715 -902 -711
rect -898 -715 -873 -711
rect -807 -715 -747 -711
rect -743 -715 -718 -711
rect -962 -721 -958 -715
rect -938 -721 -934 -715
rect -905 -721 -902 -715
rect -807 -721 -803 -715
rect -783 -721 -779 -715
rect -949 -732 -945 -725
rect -750 -721 -747 -715
rect -967 -736 -956 -732
rect -949 -735 -934 -732
rect -938 -738 -934 -735
rect -963 -744 -945 -740
rect -938 -741 -933 -738
rect -889 -741 -886 -726
rect -794 -732 -790 -725
rect -808 -736 -801 -732
rect -794 -735 -779 -732
rect -783 -738 -779 -735
rect -938 -745 -898 -741
rect -889 -744 -863 -741
rect -809 -744 -790 -740
rect -783 -741 -778 -738
rect -734 -740 -731 -726
rect -938 -752 -934 -745
rect -961 -765 -957 -756
rect -889 -760 -886 -744
rect -961 -766 -929 -765
rect -905 -766 -901 -765
rect -961 -768 -901 -766
rect -933 -769 -901 -768
rect -866 -792 -863 -744
rect -783 -745 -743 -741
rect -734 -744 -729 -740
rect -783 -752 -779 -745
rect -806 -765 -802 -756
rect -734 -760 -731 -744
rect -806 -768 -760 -765
rect -779 -769 -759 -768
rect -750 -769 -746 -765
rect -779 -770 -746 -769
rect -778 -772 -746 -770
rect -778 -773 -718 -772
rect -760 -778 -718 -773
rect -615 -792 -612 -681
rect -590 -685 -587 -681
rect -565 -683 -561 -680
rect -513 -682 -505 -678
rect -498 -681 -483 -678
rect -261 -681 -240 -677
rect -56 -673 -52 -670
rect -39 -673 -35 -663
rect -22 -666 -18 -663
rect -3 -666 1 -655
rect 101 -662 113 -661
rect -236 -677 -232 -674
rect -219 -676 -213 -674
rect -220 -677 -213 -676
rect -56 -677 -35 -673
rect 91 -663 184 -662
rect 91 -666 197 -663
rect -31 -673 -27 -670
rect -12 -671 -8 -670
rect -15 -673 -8 -671
rect -31 -674 -8 -673
rect -32 -677 -8 -674
rect 91 -672 95 -666
rect 115 -672 119 -666
rect 169 -667 197 -666
rect 169 -673 173 -667
rect 193 -673 197 -667
rect -236 -681 -213 -677
rect -590 -689 -572 -685
rect -565 -686 -560 -683
rect -513 -686 -509 -682
rect -487 -684 -483 -681
rect 104 -683 108 -676
rect -487 -686 -482 -684
rect -565 -690 -553 -686
rect -513 -690 -494 -686
rect -487 -689 -475 -686
rect -565 -697 -561 -690
rect -588 -710 -584 -701
rect -588 -713 -559 -710
rect -581 -715 -571 -713
rect -556 -780 -553 -690
rect -487 -698 -483 -689
rect -510 -711 -506 -702
rect -510 -714 -481 -711
rect -501 -716 -493 -714
rect -478 -740 -475 -689
rect 65 -687 97 -683
rect 104 -686 119 -683
rect 182 -684 186 -677
rect -117 -717 -105 -716
rect -282 -721 -222 -717
rect -218 -721 -193 -717
rect -127 -721 -67 -717
rect -63 -721 -38 -717
rect -282 -727 -278 -721
rect -258 -727 -254 -721
rect -225 -727 -222 -721
rect -127 -727 -123 -721
rect -103 -727 -99 -721
rect -269 -738 -265 -731
rect -70 -727 -67 -721
rect -550 -743 -475 -740
rect -287 -742 -276 -738
rect -269 -741 -254 -738
rect -550 -772 -546 -743
rect -258 -744 -254 -741
rect -525 -751 -514 -748
rect -283 -750 -265 -746
rect -258 -747 -253 -744
rect -209 -747 -206 -732
rect -114 -738 -110 -731
rect -128 -742 -121 -738
rect -114 -741 -99 -738
rect -103 -744 -99 -741
rect -258 -751 -218 -747
rect -209 -750 -183 -747
rect -133 -750 -110 -746
rect -103 -747 -98 -744
rect -54 -746 -51 -732
rect -532 -755 -504 -751
rect -532 -761 -528 -755
rect -508 -761 -504 -755
rect -258 -758 -254 -751
rect -519 -772 -515 -765
rect -281 -771 -277 -762
rect -209 -766 -206 -750
rect -281 -772 -249 -771
rect -225 -772 -221 -771
rect -550 -776 -526 -772
rect -519 -775 -504 -772
rect -281 -774 -221 -772
rect -253 -775 -221 -774
rect -508 -778 -504 -775
rect -556 -784 -515 -780
rect -508 -782 -480 -778
rect -508 -792 -504 -782
rect -866 -795 -612 -792
rect -531 -805 -527 -796
rect -531 -808 -502 -805
rect -520 -810 -509 -808
rect -484 -851 -480 -782
rect -186 -798 -183 -750
rect -103 -751 -63 -747
rect -54 -750 -49 -746
rect -103 -758 -99 -751
rect -126 -771 -122 -762
rect -54 -766 -51 -750
rect -126 -773 -97 -771
rect -70 -773 -66 -771
rect -126 -774 -66 -773
rect -101 -776 -66 -774
rect 65 -798 68 -687
rect 90 -691 93 -687
rect 115 -689 119 -686
rect 167 -688 175 -684
rect 182 -687 197 -684
rect 90 -695 108 -691
rect 115 -692 120 -689
rect 167 -692 171 -688
rect 193 -690 197 -687
rect 193 -692 198 -690
rect 115 -696 127 -692
rect 167 -696 186 -692
rect 193 -695 205 -692
rect 115 -703 119 -696
rect 92 -716 96 -707
rect 92 -719 121 -716
rect 99 -721 109 -719
rect 124 -786 127 -696
rect 193 -704 197 -695
rect 170 -717 174 -708
rect 170 -720 199 -717
rect 179 -722 187 -720
rect 202 -746 205 -695
rect 130 -749 205 -746
rect 130 -778 134 -749
rect 155 -757 166 -754
rect 148 -761 176 -757
rect 148 -767 152 -761
rect 172 -767 176 -761
rect 161 -778 165 -771
rect 130 -782 154 -778
rect 161 -781 176 -778
rect 172 -784 176 -781
rect 124 -790 165 -786
rect 172 -788 184 -784
rect 172 -798 176 -788
rect -186 -801 68 -798
rect 149 -811 153 -802
rect 149 -814 178 -811
rect 160 -816 171 -814
rect -1083 -855 -480 -851
rect -1902 -882 -1262 -878
<< metal2 >>
rect -666 -358 249 -354
rect -1445 -369 -1236 -365
rect -2185 -385 -1976 -381
rect -2510 -455 -2336 -451
rect -2510 -718 -2506 -455
rect -2340 -473 -2336 -455
rect -2363 -621 -2240 -617
rect -2363 -639 -2359 -621
rect -2244 -628 -2240 -621
rect -2447 -643 -2359 -639
rect -2421 -718 -2418 -683
rect -2510 -721 -2418 -718
rect -2510 -767 -2506 -721
rect -2362 -759 -2359 -643
rect -2216 -683 -2214 -679
rect -2216 -719 -2212 -683
rect -2185 -719 -2181 -385
rect -2216 -723 -2181 -719
rect -2173 -670 -2048 -667
rect -2362 -763 -2332 -759
rect -2510 -771 -2487 -767
rect -2343 -771 -2332 -767
rect -2173 -768 -2170 -670
rect -2051 -705 -2048 -670
rect -2051 -709 -2036 -705
rect -2244 -771 -2170 -768
rect -2343 -855 -2339 -771
rect -1984 -855 -1980 -385
rect -1770 -439 -1596 -435
rect -1770 -702 -1766 -439
rect -1600 -457 -1596 -439
rect -1623 -605 -1500 -601
rect -1623 -623 -1619 -605
rect -1504 -612 -1500 -605
rect -1707 -627 -1619 -623
rect -1681 -702 -1678 -667
rect -1770 -705 -1678 -702
rect -1770 -751 -1766 -705
rect -1622 -743 -1619 -627
rect -1476 -667 -1474 -663
rect -1476 -703 -1472 -667
rect -1445 -703 -1441 -369
rect -1476 -707 -1441 -703
rect -1433 -654 -1308 -651
rect -1622 -747 -1592 -743
rect -1770 -755 -1747 -751
rect -1603 -755 -1592 -751
rect -1433 -752 -1430 -654
rect -1311 -689 -1308 -654
rect -1311 -693 -1296 -689
rect -1504 -755 -1430 -752
rect -1603 -839 -1599 -755
rect -1244 -839 -1240 -369
rect -991 -428 -817 -424
rect -991 -691 -987 -428
rect -821 -446 -817 -428
rect -844 -594 -721 -590
rect -844 -612 -840 -594
rect -725 -601 -721 -594
rect -928 -616 -840 -612
rect -902 -691 -899 -656
rect -991 -694 -899 -691
rect -991 -740 -987 -694
rect -843 -732 -840 -616
rect -697 -656 -695 -652
rect -697 -692 -693 -656
rect -666 -692 -662 -358
rect -697 -696 -662 -692
rect -654 -643 -529 -640
rect -843 -736 -813 -732
rect -991 -744 -968 -740
rect -824 -744 -813 -740
rect -654 -741 -651 -643
rect -532 -678 -529 -643
rect -532 -682 -517 -678
rect -725 -744 -651 -741
rect -824 -828 -820 -744
rect -416 -828 -412 -358
rect -311 -434 -137 -430
rect -311 -697 -307 -434
rect -141 -452 -137 -434
rect -164 -600 -41 -596
rect -164 -618 -160 -600
rect -45 -607 -41 -600
rect -248 -622 -160 -618
rect -222 -697 -219 -662
rect -311 -700 -219 -697
rect -311 -746 -307 -700
rect -163 -738 -160 -622
rect 26 -649 151 -646
rect -163 -742 -133 -738
rect -311 -750 -288 -746
rect 26 -747 29 -649
rect 148 -684 151 -649
rect 148 -688 163 -684
rect -45 -750 29 -747
rect 245 -784 249 -358
rect 189 -788 249 -784
rect -824 -832 -412 -828
rect -1603 -843 -1240 -839
rect -2343 -859 -1980 -855
<< ntransistor >>
rect -2348 -529 -2346 -524
rect -2329 -529 -2327 -524
rect -2304 -529 -2302 -524
rect -2285 -529 -2283 -524
rect -1608 -513 -1606 -508
rect -1589 -513 -1587 -508
rect -1564 -513 -1562 -508
rect -1545 -513 -1543 -508
rect -829 -502 -827 -497
rect -810 -502 -808 -497
rect -785 -502 -783 -497
rect -766 -502 -764 -497
rect -149 -508 -147 -503
rect -130 -508 -128 -503
rect -105 -508 -103 -503
rect -86 -508 -84 -503
rect -2474 -695 -2472 -690
rect -2455 -695 -2453 -690
rect -2430 -695 -2428 -690
rect -2411 -695 -2409 -690
rect -2269 -691 -2267 -686
rect -2250 -691 -2248 -686
rect -2225 -691 -2223 -686
rect -2206 -691 -2204 -686
rect -1734 -679 -1732 -674
rect -1715 -679 -1713 -674
rect -1690 -679 -1688 -674
rect -1671 -679 -1669 -674
rect -1529 -675 -1527 -670
rect -1510 -675 -1508 -670
rect -1485 -675 -1483 -670
rect -1466 -675 -1464 -670
rect -2101 -733 -2098 -724
rect -2090 -733 -2087 -724
rect -955 -668 -953 -663
rect -936 -668 -934 -663
rect -911 -668 -909 -663
rect -892 -668 -890 -663
rect -750 -664 -748 -659
rect -731 -664 -729 -659
rect -706 -664 -704 -659
rect -687 -664 -685 -659
rect -1361 -717 -1358 -708
rect -1350 -717 -1347 -708
rect -582 -706 -579 -697
rect -571 -706 -568 -697
rect -275 -674 -273 -669
rect -256 -674 -254 -669
rect -231 -674 -229 -669
rect -212 -674 -210 -669
rect -70 -670 -68 -665
rect -51 -670 -49 -665
rect -26 -670 -24 -665
rect -7 -670 -5 -665
rect -504 -707 -501 -698
rect -493 -707 -490 -698
rect -1283 -718 -1280 -709
rect -1272 -718 -1269 -709
rect 98 -712 101 -703
rect 109 -712 112 -703
rect 176 -713 179 -704
rect 187 -713 190 -704
rect -2023 -734 -2020 -725
rect -2012 -734 -2009 -725
rect -2474 -788 -2471 -779
rect -2463 -788 -2460 -779
rect -1734 -772 -1731 -763
rect -1723 -772 -1720 -763
rect -2416 -792 -2413 -787
rect -2319 -788 -2316 -779
rect -2308 -788 -2305 -779
rect -1676 -776 -1673 -771
rect -1579 -772 -1576 -763
rect -1568 -772 -1565 -763
rect -955 -761 -952 -752
rect -944 -761 -941 -752
rect -897 -765 -894 -760
rect -800 -761 -797 -752
rect -789 -761 -786 -752
rect -742 -765 -739 -760
rect -1521 -776 -1518 -771
rect -275 -767 -272 -758
rect -264 -767 -261 -758
rect -2261 -792 -2258 -787
rect -217 -771 -214 -766
rect -120 -767 -117 -758
rect -109 -767 -106 -758
rect -62 -771 -59 -766
rect -525 -801 -522 -792
rect -514 -801 -511 -792
rect -1304 -812 -1301 -803
rect -1293 -812 -1290 -803
rect 155 -807 158 -798
rect 166 -807 169 -798
rect -2044 -828 -2041 -819
rect -2033 -828 -2030 -819
<< ptransistor >>
rect -2348 -498 -2346 -493
rect -2329 -498 -2327 -493
rect -2304 -498 -2302 -493
rect -2285 -498 -2283 -493
rect -1608 -482 -1606 -477
rect -1589 -482 -1587 -477
rect -1564 -482 -1562 -477
rect -1545 -482 -1543 -477
rect -829 -471 -827 -466
rect -810 -471 -808 -466
rect -785 -471 -783 -466
rect -766 -471 -764 -466
rect -149 -477 -147 -472
rect -130 -477 -128 -472
rect -105 -477 -103 -472
rect -86 -477 -84 -472
rect -2474 -664 -2472 -659
rect -2455 -664 -2453 -659
rect -2430 -664 -2428 -659
rect -2411 -664 -2409 -659
rect -2269 -660 -2267 -655
rect -2250 -660 -2248 -655
rect -2225 -660 -2223 -655
rect -2206 -660 -2204 -655
rect -2101 -700 -2098 -693
rect -2090 -700 -2087 -693
rect -1734 -648 -1732 -643
rect -1715 -648 -1713 -643
rect -1690 -648 -1688 -643
rect -1671 -648 -1669 -643
rect -1529 -644 -1527 -639
rect -1510 -644 -1508 -639
rect -1485 -644 -1483 -639
rect -1466 -644 -1464 -639
rect -1361 -684 -1358 -677
rect -1350 -684 -1347 -677
rect -2023 -701 -2020 -694
rect -2012 -701 -2009 -694
rect -1283 -685 -1280 -678
rect -1272 -685 -1269 -678
rect -955 -637 -953 -632
rect -936 -637 -934 -632
rect -911 -637 -909 -632
rect -892 -637 -890 -632
rect -750 -633 -748 -628
rect -731 -633 -729 -628
rect -706 -633 -704 -628
rect -687 -633 -685 -628
rect -582 -673 -579 -666
rect -571 -673 -568 -666
rect -504 -674 -501 -667
rect -493 -674 -490 -667
rect -275 -643 -273 -638
rect -256 -643 -254 -638
rect -231 -643 -229 -638
rect -212 -643 -210 -638
rect -70 -639 -68 -634
rect -51 -639 -49 -634
rect -26 -639 -24 -634
rect -7 -639 -5 -634
rect 98 -679 101 -672
rect 109 -679 112 -672
rect 176 -680 179 -673
rect 187 -680 190 -673
rect -955 -728 -952 -721
rect -944 -728 -941 -721
rect -897 -726 -894 -721
rect -1734 -739 -1731 -732
rect -1723 -739 -1720 -732
rect -1676 -737 -1673 -732
rect -2474 -755 -2471 -748
rect -2463 -755 -2460 -748
rect -2416 -753 -2413 -748
rect -2319 -755 -2316 -748
rect -2308 -755 -2305 -748
rect -2261 -753 -2258 -748
rect -1579 -739 -1576 -732
rect -1568 -739 -1565 -732
rect -1521 -737 -1518 -732
rect -800 -728 -797 -721
rect -789 -728 -786 -721
rect -742 -726 -739 -721
rect -275 -734 -272 -727
rect -264 -734 -261 -727
rect -217 -732 -214 -727
rect -120 -734 -117 -727
rect -109 -734 -106 -727
rect -62 -732 -59 -727
rect -525 -768 -522 -761
rect -514 -768 -511 -761
rect -1304 -779 -1301 -772
rect -1293 -779 -1290 -772
rect -2044 -795 -2041 -788
rect -2033 -795 -2030 -788
rect 155 -774 158 -767
rect 166 -774 169 -767
<< polycontact >>
rect -2307 -514 -2303 -510
rect -2288 -514 -2284 -510
rect -2278 -514 -2274 -510
rect -1567 -498 -1563 -494
rect -1548 -498 -1544 -494
rect -1538 -498 -1534 -494
rect -788 -487 -784 -483
rect -769 -487 -765 -483
rect -759 -487 -755 -483
rect -108 -493 -104 -489
rect -89 -493 -85 -489
rect -79 -493 -75 -489
rect -2433 -680 -2429 -676
rect -2414 -681 -2410 -677
rect -2404 -680 -2400 -676
rect -2228 -676 -2224 -672
rect -2209 -676 -2205 -672
rect -2199 -676 -2195 -672
rect -1693 -664 -1689 -660
rect -1674 -665 -1670 -661
rect -1664 -664 -1660 -660
rect -1488 -660 -1484 -656
rect -1469 -660 -1465 -656
rect -1459 -660 -1455 -656
rect -1362 -692 -1358 -688
rect -2102 -708 -2098 -704
rect -2024 -709 -2020 -705
rect -2091 -716 -2087 -712
rect -914 -653 -910 -649
rect -895 -654 -891 -650
rect -885 -653 -881 -649
rect -709 -649 -705 -645
rect -690 -649 -686 -645
rect -680 -649 -676 -645
rect -583 -681 -579 -677
rect -1284 -693 -1280 -689
rect -1351 -700 -1347 -696
rect -2013 -717 -2009 -713
rect -505 -682 -501 -678
rect -572 -689 -568 -685
rect -1273 -701 -1269 -697
rect -494 -690 -490 -686
rect -234 -659 -230 -655
rect -215 -660 -211 -656
rect -205 -659 -201 -655
rect -29 -655 -25 -651
rect -10 -655 -6 -651
rect 0 -655 4 -651
rect 97 -687 101 -683
rect 175 -688 179 -684
rect 108 -695 112 -691
rect 186 -696 190 -692
rect -1735 -747 -1731 -743
rect -2475 -763 -2471 -759
rect -2464 -771 -2460 -767
rect -2320 -763 -2316 -759
rect -2417 -772 -2413 -768
rect -2309 -771 -2305 -767
rect -1724 -755 -1720 -751
rect -956 -736 -952 -732
rect -1580 -747 -1576 -743
rect -1677 -756 -1673 -752
rect -2262 -772 -2258 -768
rect -1569 -755 -1565 -751
rect -945 -744 -941 -740
rect -801 -736 -797 -732
rect -898 -745 -894 -741
rect -1522 -756 -1518 -752
rect -790 -744 -786 -740
rect -743 -745 -739 -741
rect -276 -742 -272 -738
rect -265 -750 -261 -746
rect -121 -742 -117 -738
rect -218 -751 -214 -747
rect -110 -750 -106 -746
rect -63 -751 -59 -747
rect -526 -776 -522 -772
rect -1305 -787 -1301 -783
rect -2045 -803 -2041 -799
rect -1294 -795 -1290 -791
rect -515 -784 -511 -780
rect 154 -782 158 -778
rect 165 -790 169 -786
rect -2034 -811 -2030 -807
<< ndcontact >>
rect -2353 -529 -2349 -525
rect -2344 -529 -2340 -525
rect -2334 -529 -2330 -525
rect -2325 -529 -2321 -525
rect -2309 -529 -2305 -525
rect -2300 -529 -2296 -525
rect -2290 -529 -2286 -525
rect -2281 -529 -2277 -525
rect -1613 -513 -1609 -509
rect -1604 -513 -1600 -509
rect -1594 -513 -1590 -509
rect -1585 -513 -1581 -509
rect -1569 -513 -1565 -509
rect -1560 -513 -1556 -509
rect -1550 -513 -1546 -509
rect -1541 -513 -1537 -509
rect -834 -502 -830 -498
rect -825 -502 -821 -498
rect -815 -502 -811 -498
rect -806 -502 -802 -498
rect -790 -502 -786 -498
rect -781 -502 -777 -498
rect -771 -502 -767 -498
rect -762 -502 -758 -498
rect -154 -508 -150 -504
rect -145 -508 -141 -504
rect -135 -508 -131 -504
rect -126 -508 -122 -504
rect -110 -508 -106 -504
rect -101 -508 -97 -504
rect -91 -508 -87 -504
rect -82 -508 -78 -504
rect -2479 -695 -2475 -691
rect -2470 -695 -2466 -691
rect -2460 -695 -2456 -691
rect -2451 -695 -2447 -691
rect -2435 -695 -2431 -691
rect -2426 -695 -2422 -691
rect -2416 -695 -2412 -691
rect -2407 -695 -2403 -691
rect -2274 -691 -2270 -687
rect -2265 -691 -2261 -687
rect -2255 -691 -2251 -687
rect -2246 -691 -2242 -687
rect -2230 -691 -2226 -687
rect -2221 -691 -2217 -687
rect -2211 -691 -2207 -687
rect -2202 -691 -2198 -687
rect -1739 -679 -1735 -675
rect -1730 -679 -1726 -675
rect -1720 -679 -1716 -675
rect -1711 -679 -1707 -675
rect -1695 -679 -1691 -675
rect -1686 -679 -1682 -675
rect -1676 -679 -1672 -675
rect -1667 -679 -1663 -675
rect -1534 -675 -1530 -671
rect -1525 -675 -1521 -671
rect -1515 -675 -1511 -671
rect -1506 -675 -1502 -671
rect -1490 -675 -1486 -671
rect -1481 -675 -1477 -671
rect -1471 -675 -1467 -671
rect -1462 -675 -1458 -671
rect -2107 -728 -2103 -724
rect -2084 -728 -2080 -724
rect -960 -668 -956 -664
rect -951 -668 -947 -664
rect -941 -668 -937 -664
rect -932 -668 -928 -664
rect -916 -668 -912 -664
rect -907 -668 -903 -664
rect -897 -668 -893 -664
rect -888 -668 -884 -664
rect -755 -664 -751 -660
rect -746 -664 -742 -660
rect -736 -664 -732 -660
rect -727 -664 -723 -660
rect -711 -664 -707 -660
rect -702 -664 -698 -660
rect -692 -664 -688 -660
rect -683 -664 -679 -660
rect -1367 -712 -1363 -708
rect -1344 -712 -1340 -708
rect -588 -701 -584 -697
rect -565 -701 -561 -697
rect -280 -674 -276 -670
rect -271 -674 -267 -670
rect -261 -674 -257 -670
rect -252 -674 -248 -670
rect -236 -674 -232 -670
rect -227 -674 -223 -670
rect -217 -674 -213 -670
rect -208 -674 -204 -670
rect -75 -670 -71 -666
rect -66 -670 -62 -666
rect -56 -670 -52 -666
rect -47 -670 -43 -666
rect -31 -670 -27 -666
rect -22 -670 -18 -666
rect -12 -670 -8 -666
rect -3 -670 1 -666
rect -510 -702 -506 -698
rect -487 -702 -483 -698
rect 92 -707 96 -703
rect -1289 -713 -1285 -709
rect -1266 -713 -1262 -709
rect 115 -707 119 -703
rect 170 -708 174 -704
rect 193 -708 197 -704
rect -2029 -729 -2025 -725
rect -2006 -729 -2002 -725
rect -2480 -783 -2476 -779
rect -2457 -783 -2453 -779
rect -1740 -767 -1736 -763
rect -1717 -767 -1713 -763
rect -1585 -767 -1581 -763
rect -2325 -783 -2321 -779
rect -2424 -792 -2419 -787
rect -2409 -792 -2405 -787
rect -2302 -783 -2298 -779
rect -1684 -776 -1679 -771
rect -1669 -776 -1665 -771
rect -1562 -767 -1558 -763
rect -961 -756 -957 -752
rect -938 -756 -934 -752
rect -806 -756 -802 -752
rect -905 -765 -900 -760
rect -890 -765 -886 -760
rect -783 -756 -779 -752
rect -750 -765 -745 -760
rect -735 -765 -731 -760
rect -1529 -776 -1524 -771
rect -1514 -776 -1510 -771
rect -281 -762 -277 -758
rect -258 -762 -254 -758
rect -126 -762 -122 -758
rect -2269 -792 -2264 -787
rect -2254 -792 -2250 -787
rect -225 -771 -220 -766
rect -210 -771 -206 -766
rect -103 -762 -99 -758
rect -70 -771 -65 -766
rect -55 -771 -51 -766
rect -531 -796 -527 -792
rect -508 -796 -504 -792
rect -1310 -807 -1306 -803
rect -1287 -807 -1283 -803
rect 149 -802 153 -798
rect 172 -802 176 -798
rect -2050 -823 -2046 -819
rect -2027 -823 -2023 -819
<< pdcontact >>
rect -2353 -498 -2349 -494
rect -2344 -498 -2340 -494
rect -2334 -498 -2330 -494
rect -2325 -498 -2321 -494
rect -2309 -498 -2305 -494
rect -2300 -498 -2296 -494
rect -2290 -498 -2286 -494
rect -2281 -498 -2277 -494
rect -1613 -482 -1609 -478
rect -1604 -482 -1600 -478
rect -1594 -482 -1590 -478
rect -1585 -482 -1581 -478
rect -1569 -482 -1565 -478
rect -1560 -482 -1556 -478
rect -1550 -482 -1546 -478
rect -1541 -482 -1537 -478
rect -834 -471 -830 -467
rect -825 -471 -821 -467
rect -815 -471 -811 -467
rect -806 -471 -802 -467
rect -790 -471 -786 -467
rect -781 -471 -777 -467
rect -771 -471 -767 -467
rect -762 -471 -758 -467
rect -154 -477 -150 -473
rect -145 -477 -141 -473
rect -135 -477 -131 -473
rect -126 -477 -122 -473
rect -110 -477 -106 -473
rect -101 -477 -97 -473
rect -91 -477 -87 -473
rect -82 -477 -78 -473
rect -2479 -664 -2475 -660
rect -2470 -664 -2466 -660
rect -2460 -664 -2456 -660
rect -2451 -664 -2447 -660
rect -2435 -664 -2431 -660
rect -2426 -664 -2422 -660
rect -2416 -664 -2412 -660
rect -2407 -664 -2403 -660
rect -2274 -660 -2270 -656
rect -2265 -660 -2261 -656
rect -2255 -660 -2251 -656
rect -2246 -660 -2242 -656
rect -2230 -660 -2226 -656
rect -2221 -660 -2217 -656
rect -2211 -660 -2207 -656
rect -2202 -660 -2198 -656
rect -2108 -697 -2104 -693
rect -2095 -697 -2091 -693
rect -2084 -697 -2080 -693
rect -1739 -648 -1735 -644
rect -1730 -648 -1726 -644
rect -1720 -648 -1716 -644
rect -1711 -648 -1707 -644
rect -1695 -648 -1691 -644
rect -1686 -648 -1682 -644
rect -1676 -648 -1672 -644
rect -1667 -648 -1663 -644
rect -1534 -644 -1530 -640
rect -1525 -644 -1521 -640
rect -1515 -644 -1511 -640
rect -1506 -644 -1502 -640
rect -1490 -644 -1486 -640
rect -1481 -644 -1477 -640
rect -1471 -644 -1467 -640
rect -1462 -644 -1458 -640
rect -1368 -681 -1364 -677
rect -1355 -681 -1351 -677
rect -1344 -681 -1340 -677
rect -1290 -682 -1286 -678
rect -2030 -698 -2026 -694
rect -2017 -698 -2013 -694
rect -2006 -698 -2002 -694
rect -1277 -682 -1273 -678
rect -1266 -682 -1262 -678
rect -960 -637 -956 -633
rect -951 -637 -947 -633
rect -941 -637 -937 -633
rect -932 -637 -928 -633
rect -916 -637 -912 -633
rect -907 -637 -903 -633
rect -897 -637 -893 -633
rect -888 -637 -884 -633
rect -755 -633 -751 -629
rect -746 -633 -742 -629
rect -736 -633 -732 -629
rect -727 -633 -723 -629
rect -711 -633 -707 -629
rect -702 -633 -698 -629
rect -692 -633 -688 -629
rect -683 -633 -679 -629
rect -589 -670 -585 -666
rect -576 -670 -572 -666
rect -565 -670 -561 -666
rect -511 -671 -507 -667
rect -498 -671 -494 -667
rect -487 -671 -483 -667
rect -280 -643 -276 -639
rect -271 -643 -267 -639
rect -261 -643 -257 -639
rect -252 -643 -248 -639
rect -236 -643 -232 -639
rect -227 -643 -223 -639
rect -217 -643 -213 -639
rect -208 -643 -204 -639
rect -75 -639 -71 -635
rect -66 -639 -62 -635
rect -56 -639 -52 -635
rect -47 -639 -43 -635
rect -31 -639 -27 -635
rect -22 -639 -18 -635
rect -12 -639 -8 -635
rect -3 -639 1 -635
rect 91 -676 95 -672
rect 104 -676 108 -672
rect 115 -676 119 -672
rect 169 -677 173 -673
rect 182 -677 186 -673
rect 193 -677 197 -673
rect -962 -725 -958 -721
rect -949 -725 -945 -721
rect -938 -725 -934 -721
rect -905 -726 -901 -721
rect -890 -726 -886 -721
rect -807 -725 -803 -721
rect -1741 -736 -1737 -732
rect -1728 -736 -1724 -732
rect -1717 -736 -1713 -732
rect -1684 -737 -1680 -732
rect -1669 -737 -1665 -732
rect -1586 -736 -1582 -732
rect -2481 -752 -2477 -748
rect -2468 -752 -2464 -748
rect -2457 -752 -2453 -748
rect -2424 -753 -2420 -748
rect -2409 -753 -2405 -748
rect -2326 -752 -2322 -748
rect -2313 -752 -2309 -748
rect -2302 -752 -2298 -748
rect -2269 -753 -2265 -748
rect -2254 -753 -2250 -748
rect -1573 -736 -1569 -732
rect -1562 -736 -1558 -732
rect -1529 -737 -1525 -732
rect -1514 -737 -1510 -732
rect -794 -725 -790 -721
rect -783 -725 -779 -721
rect -750 -726 -746 -721
rect -735 -726 -731 -721
rect -282 -731 -278 -727
rect -269 -731 -265 -727
rect -258 -731 -254 -727
rect -225 -732 -221 -727
rect -210 -732 -206 -727
rect -127 -731 -123 -727
rect -114 -731 -110 -727
rect -103 -731 -99 -727
rect -70 -732 -66 -727
rect -55 -732 -51 -727
rect -532 -765 -528 -761
rect -519 -765 -515 -761
rect -508 -765 -504 -761
rect -1311 -776 -1307 -772
rect -1298 -776 -1294 -772
rect -1287 -776 -1283 -772
rect -2051 -792 -2047 -788
rect -2038 -792 -2034 -788
rect -2027 -792 -2023 -788
rect 148 -771 152 -767
rect 161 -771 165 -767
rect 172 -771 176 -767
<< m2contact >>
rect -1236 -369 -1232 -365
rect -1976 -385 -1972 -381
rect -2340 -477 -2336 -473
rect -2244 -632 -2240 -628
rect -2451 -643 -2447 -639
rect -2418 -687 -2414 -683
rect -2214 -683 -2210 -679
rect -2487 -771 -2482 -767
rect -2332 -763 -2327 -759
rect -2332 -771 -2328 -767
rect -2248 -771 -2244 -767
rect -2036 -709 -2032 -705
rect -1600 -461 -1596 -457
rect -1504 -616 -1500 -612
rect -1711 -627 -1707 -623
rect -1678 -671 -1674 -667
rect -1474 -667 -1470 -663
rect -1747 -755 -1742 -751
rect -1592 -747 -1587 -743
rect -1592 -755 -1588 -751
rect -1508 -755 -1504 -751
rect -1296 -693 -1292 -689
rect -821 -450 -817 -446
rect -141 -456 -137 -452
rect -725 -605 -721 -601
rect -932 -616 -928 -612
rect -899 -660 -895 -656
rect -45 -611 -41 -607
rect -695 -656 -691 -652
rect -252 -622 -248 -618
rect -219 -666 -215 -662
rect -968 -744 -963 -740
rect -813 -736 -808 -732
rect -813 -744 -809 -740
rect -729 -744 -725 -740
rect -517 -682 -513 -678
rect -288 -750 -283 -746
rect -133 -742 -128 -738
rect -49 -750 -45 -746
rect 163 -688 167 -684
rect 184 -788 189 -784
<< nsubstratencontact >>
rect -902 -715 -898 -711
rect -747 -715 -743 -711
rect -222 -721 -218 -717
rect -67 -721 -63 -717
rect -1681 -726 -1677 -722
rect -1526 -726 -1522 -722
rect -2421 -742 -2417 -738
rect -2266 -742 -2262 -738
<< labels >>
rlabel metal1 -778 -506 -778 -506 1 gnd
rlabel metal1 -779 -453 -779 -453 1 vdd
rlabel metal1 -770 -485 -770 -485 1 M
rlabel metal1 -907 -673 -907 -673 1 gnd
rlabel metal1 -908 -619 -908 -619 1 vdd
rlabel metal1 -924 -713 -924 -713 1 vdd
rlabel metal1 -924 -768 -924 -768 1 gnd
rlabel metal1 -698 -614 -698 -614 1 vdd
rlabel metal1 -699 -669 -699 -669 1 gnd
rlabel metal1 -795 -484 -795 -484 1 B1
rlabel metal1 -923 -651 -923 -651 1 A1
rlabel metal1 -964 -734 -964 -734 1 A1
rlabel metal1 -739 -610 -739 -610 1 S1
rlabel metal1 -768 -712 -768 -712 1 vdd
rlabel metal1 -764 -769 -763 -768 1 gnd
rlabel metal1 -553 -658 -553 -658 1 vdd
rlabel metal1 -575 -714 -575 -714 1 gnd
rlabel metal1 -497 -715 -497 -715 1 gnd
rlabel metal1 -516 -807 -516 -807 1 gnd
rlabel metal1 -520 -750 -520 -750 1 vdd
rlabel metal1 -495 -779 -495 -779 1 C2
rlabel metal1 -1557 -517 -1557 -517 1 gnd
rlabel metal1 -1558 -464 -1558 -464 1 vdd
rlabel metal1 -1549 -496 -1549 -496 1 M
rlabel metal1 -1686 -684 -1686 -684 1 gnd
rlabel metal1 -1687 -630 -1687 -630 1 vdd
rlabel metal1 -1703 -724 -1703 -724 1 vdd
rlabel metal1 -1703 -779 -1703 -779 1 gnd
rlabel metal1 -1477 -625 -1477 -625 1 vdd
rlabel metal1 -1478 -680 -1478 -680 1 gnd
rlabel metal1 -1547 -723 -1547 -723 1 vdd
rlabel metal1 -1543 -780 -1542 -779 1 gnd
rlabel metal1 -1332 -669 -1332 -669 1 vdd
rlabel metal1 -1354 -725 -1354 -725 1 gnd
rlabel metal1 -1276 -726 -1276 -726 1 gnd
rlabel metal1 -1295 -818 -1295 -818 1 gnd
rlabel metal1 -1299 -761 -1299 -761 1 vdd
rlabel metal1 -1575 -495 -1575 -495 1 B2
rlabel metal1 -1701 -661 -1701 -661 1 A2
rlabel metal1 -1743 -745 -1743 -745 1 A2
rlabel metal1 -1518 -622 -1518 -622 1 S2
rlabel metal1 -1274 -790 -1274 -790 1 C3
rlabel metal1 -2297 -533 -2297 -533 1 gnd
rlabel metal1 -2298 -480 -2298 -480 1 vdd
rlabel metal1 -2289 -512 -2289 -512 1 M
rlabel metal1 -2426 -700 -2426 -700 1 gnd
rlabel metal1 -2427 -646 -2427 -646 1 vdd
rlabel metal1 -2443 -740 -2443 -740 1 vdd
rlabel metal1 -2443 -795 -2443 -795 1 gnd
rlabel metal1 -2217 -641 -2217 -641 1 vdd
rlabel metal1 -2218 -696 -2218 -696 1 gnd
rlabel metal1 -2287 -739 -2287 -739 1 vdd
rlabel metal1 -2283 -796 -2282 -795 1 gnd
rlabel metal1 -2072 -685 -2072 -685 1 vdd
rlabel metal1 -2094 -741 -2094 -741 1 gnd
rlabel metal1 -2016 -742 -2016 -742 1 gnd
rlabel metal1 -2035 -834 -2035 -834 1 gnd
rlabel metal1 -2039 -777 -2039 -777 1 vdd
rlabel metal1 -2314 -512 -2314 -512 1 B3
rlabel metal1 -2440 -677 -2440 -677 1 A3
rlabel metal1 -2483 -761 -2483 -761 1 A3
rlabel metal1 -2257 -637 -2257 -637 1 S3
rlabel metal1 -2012 -807 -2012 -807 1 carry
rlabel metal1 -98 -512 -98 -512 1 gnd
rlabel metal1 -99 -459 -99 -459 1 vdd
rlabel metal1 -115 -491 -115 -491 1 B0
rlabel metal1 -90 -491 -90 -491 1 M
rlabel metal1 -227 -679 -227 -679 1 gnd
rlabel metal1 -241 -657 -241 -657 1 A0
rlabel metal1 -228 -625 -228 -625 1 vdd
rlabel metal1 -244 -719 -244 -719 1 vdd
rlabel metal1 -244 -774 -244 -774 1 gnd
rlabel metal1 -283 -740 -283 -740 1 A0
rlabel metal1 -18 -620 -18 -620 1 vdd
rlabel metal1 -19 -675 -19 -675 1 gnd
rlabel metal1 -12 -653 -12 -653 1 M
rlabel metal1 -60 -616 -60 -616 1 S0
rlabel metal1 -90 -774 -90 -774 1 gnd
rlabel metal1 -87 -719 -87 -719 1 vdd
rlabel metal1 -128 -748 -128 -748 1 M
rlabel metal1 137 -664 137 -664 1 vdd
rlabel metal1 102 -718 102 -718 1 gnd
rlabel metal1 183 -720 183 -720 1 gnd
rlabel metal1 161 -756 162 -755 1 vdd
rlabel metal1 166 -814 166 -814 1 gnd
rlabel m2contact 185 -786 185 -786 1 C1
<< end >>
