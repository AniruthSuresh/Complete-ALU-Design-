magic
tech scmos
timestamp 1701530711
<< nwell >>
rect 2981 633 3061 656
rect 3721 649 3801 672
rect 4500 660 4580 683
rect 5180 654 5260 677
rect 2855 467 2935 490
rect 3060 471 3140 494
rect 3595 483 3675 506
rect 3800 487 3880 510
rect 4374 494 4454 517
rect 4579 498 4659 521
rect 5054 488 5134 511
rect 5259 492 5339 515
rect 3963 453 4001 469
rect 1253 429 1291 445
rect 1331 428 1369 444
rect 3223 437 3261 453
rect 4041 452 4079 468
rect 4742 464 4780 480
rect 4820 463 4858 479
rect 5422 458 5460 474
rect 5500 457 5538 473
rect 3301 436 3339 452
rect 3590 398 3628 414
rect 1417 369 1455 385
rect 1469 367 1510 385
rect 1528 371 1566 387
rect 1580 369 1621 387
rect 1644 371 1682 387
rect 1696 369 1737 387
rect 1764 372 1802 388
rect 1816 370 1857 388
rect 1946 373 1984 389
rect 1998 371 2039 389
rect 2057 375 2095 391
rect 2109 373 2150 391
rect 2173 375 2211 391
rect 2225 373 2266 391
rect 2293 376 2331 392
rect 2345 374 2386 392
rect 2850 382 2888 398
rect 2902 380 2943 398
rect 3005 382 3043 398
rect 3057 380 3098 398
rect 3642 396 3683 414
rect 3745 398 3783 414
rect 3797 396 3838 414
rect 4369 409 4407 425
rect 4421 407 4462 425
rect 4524 409 4562 425
rect 4576 407 4617 425
rect 5049 403 5087 419
rect 5101 401 5142 419
rect 5204 403 5242 419
rect 5256 401 5297 419
rect 4020 358 4058 374
rect 4799 369 4837 385
rect 5479 363 5517 379
rect 1076 319 1114 335
rect 1128 317 1169 335
rect 1310 334 1348 350
rect 3280 342 3318 358
rect 971 223 1012 241
rect 1078 236 1116 252
rect 1130 234 1171 252
rect 1420 167 1458 183
rect 1472 165 1513 183
rect 1531 169 1569 185
rect 1583 167 1624 185
rect 1647 169 1685 185
rect 1699 167 1740 185
rect 1767 170 1805 186
rect 1819 168 1860 186
rect 1949 171 1987 187
rect 2001 169 2042 187
rect 2060 173 2098 189
rect 2112 171 2153 189
rect 2176 173 2214 189
rect 2228 171 2269 189
rect 2296 174 2334 190
rect 2348 172 2389 190
rect 972 126 1013 144
rect 1076 136 1114 152
rect 1128 134 1169 152
rect 1077 47 1115 63
rect 1129 45 1170 63
rect 1445 -10 1483 6
rect 1497 -12 1538 6
rect 1556 -8 1594 8
rect 1608 -10 1649 8
rect 1672 -8 1710 8
rect 1724 -10 1765 8
rect 1792 -7 1830 9
rect 1844 -9 1885 9
rect 1974 -6 2012 10
rect 2026 -8 2067 10
rect 2085 -4 2123 12
rect 2137 -6 2178 12
rect 2201 -4 2239 12
rect 2253 -6 2294 12
rect 2321 -3 2359 13
rect 2373 -5 2414 13
rect 3580 6 3618 22
rect 3658 5 3696 21
rect 3637 -89 3675 -73
rect 3798 -121 3836 -105
rect 3876 -122 3914 -106
rect 1712 -151 1750 -135
rect 1764 -153 1805 -135
rect 1830 -152 1868 -136
rect 1882 -154 1923 -136
rect 1963 -152 2001 -136
rect 2015 -154 2056 -136
rect 2082 -153 2120 -137
rect 2134 -155 2175 -137
rect 4086 -160 4127 -142
rect 3855 -216 3893 -200
rect 3593 -270 3631 -254
rect 3671 -271 3709 -255
rect 3650 -365 3688 -349
rect 2819 -604 2860 -586
rect 2984 -604 3025 -586
rect 3161 -603 3202 -585
rect 3336 -604 3377 -586
rect 3734 -649 3775 -631
rect 3824 -664 3904 -641
rect 3982 -650 4023 -632
rect 4225 -641 4266 -623
rect 4072 -665 4152 -642
rect 4315 -656 4395 -633
rect 4494 -636 4535 -618
rect 4584 -651 4664 -628
rect 2870 -721 2908 -705
rect 2922 -723 2963 -705
rect 3041 -716 3079 -700
rect 3093 -718 3134 -700
rect 3234 -720 3272 -704
rect 3286 -722 3327 -704
rect 3415 -716 3453 -700
rect 3467 -718 3508 -700
rect 4073 -777 4111 -761
rect 4125 -779 4166 -761
rect 4293 -797 4331 -781
rect 4345 -799 4386 -781
rect 4449 -789 4487 -773
rect 4501 -791 4542 -773
rect 3002 -860 3040 -844
rect 3054 -862 3095 -844
rect 3852 -892 3890 -876
rect 3904 -894 3945 -876
rect 5003 -1014 5041 -998
rect 5055 -1016 5096 -998
rect 5220 -1015 5258 -999
rect 5272 -1017 5313 -999
rect 3006 -1058 3044 -1042
rect 3058 -1060 3099 -1042
rect 4193 -1061 4231 -1045
rect 3865 -1078 3903 -1062
rect 3917 -1080 3958 -1062
rect 4245 -1063 4286 -1045
rect 2844 -1235 2885 -1217
rect 3009 -1235 3050 -1217
rect 3186 -1234 3227 -1216
rect 3361 -1235 3402 -1217
rect 2895 -1352 2933 -1336
rect 2947 -1354 2988 -1336
rect 3066 -1347 3104 -1331
rect 3118 -1349 3159 -1331
rect 3259 -1351 3297 -1335
rect 3311 -1353 3352 -1335
rect 3440 -1347 3478 -1331
rect 3492 -1349 3533 -1331
rect 3652 -1548 3690 -1532
rect 3730 -1549 3768 -1533
rect 3709 -1643 3747 -1627
rect 3997 -1658 4035 -1642
rect 4075 -1659 4113 -1643
rect 4548 -1647 4589 -1629
rect 4054 -1753 4092 -1737
rect 3662 -1792 3700 -1776
rect 3740 -1793 3778 -1777
rect 3719 -1887 3757 -1871
<< polysilicon >>
rect 3035 697 3039 986
rect 3776 708 3780 986
rect 4555 726 4559 986
rect 4555 722 4613 726
rect 3776 704 3860 708
rect 3035 693 3117 697
rect 2973 676 3009 678
rect 2973 599 2975 676
rect 2988 647 2990 649
rect 3007 647 3009 676
rect 3035 664 3039 693
rect 3032 647 3034 649
rect 3051 647 3053 649
rect 2988 630 2990 642
rect 3007 640 3009 642
rect 3032 630 3034 642
rect 3051 630 3053 642
rect 2988 628 3009 630
rect 2988 616 2990 619
rect 3007 616 3009 628
rect 3033 626 3034 630
rect 3052 626 3053 630
rect 3062 627 3068 629
rect 3032 616 3034 626
rect 3051 616 3053 626
rect 2988 599 2990 611
rect 3007 603 3009 611
rect 3032 609 3034 611
rect 3051 603 3053 611
rect 3007 601 3053 603
rect 3066 599 3068 627
rect 2973 597 3068 599
rect 3113 567 3117 693
rect 3713 692 3749 694
rect 3713 615 3715 692
rect 3728 663 3730 665
rect 3747 663 3749 692
rect 3776 680 3780 704
rect 3772 663 3774 665
rect 3791 663 3793 665
rect 3728 646 3730 658
rect 3747 656 3749 658
rect 3772 646 3774 658
rect 3791 646 3793 658
rect 3728 644 3749 646
rect 3728 632 3730 635
rect 3747 632 3749 644
rect 3773 642 3774 646
rect 3792 642 3793 646
rect 3802 643 3808 645
rect 3772 632 3774 642
rect 3791 632 3793 642
rect 3728 615 3730 627
rect 3747 619 3749 627
rect 3772 625 3774 627
rect 3791 619 3793 627
rect 3747 617 3793 619
rect 3806 615 3808 643
rect 3713 613 3808 615
rect 3856 590 3860 704
rect 4492 703 4528 705
rect 4492 626 4494 703
rect 4507 674 4509 676
rect 4526 674 4528 703
rect 4555 691 4559 722
rect 4551 674 4553 676
rect 4570 674 4572 676
rect 4507 657 4509 669
rect 4526 667 4528 669
rect 4551 657 4553 669
rect 4570 657 4572 669
rect 4507 655 4528 657
rect 4507 643 4509 646
rect 4526 643 4528 655
rect 4552 653 4553 657
rect 4571 653 4572 657
rect 4581 654 4587 656
rect 4551 643 4553 653
rect 4570 643 4572 653
rect 4507 626 4509 638
rect 4526 630 4528 638
rect 4551 636 4553 638
rect 4570 630 4572 638
rect 4526 628 4572 630
rect 4585 626 4587 654
rect 4492 624 4587 626
rect 3651 589 3860 590
rect 3651 586 4024 589
rect 2916 563 3278 567
rect 2847 510 2883 512
rect 1079 483 1301 487
rect 1079 350 1083 483
rect 1297 451 1301 483
rect 1265 439 1268 443
rect 1276 439 1279 443
rect 1265 428 1268 432
rect 1265 408 1268 424
rect 1276 420 1279 432
rect 1276 408 1279 416
rect 1265 396 1268 399
rect 1276 396 1279 399
rect 1275 389 1276 392
rect 981 346 1122 350
rect 981 274 985 346
rect 1118 341 1122 346
rect 1088 329 1091 333
rect 1099 329 1102 333
rect 1146 329 1149 332
rect 1088 318 1091 322
rect 1088 298 1091 314
rect 1099 310 1102 322
rect 1146 309 1149 324
rect 1099 298 1102 306
rect 1146 290 1149 305
rect 1088 286 1091 289
rect 1099 286 1102 289
rect 1146 282 1149 285
rect 1271 280 1276 389
rect 1316 382 1320 443
rect 1343 438 1346 442
rect 1354 438 1357 442
rect 2847 433 2849 510
rect 2862 481 2864 483
rect 2881 481 2883 510
rect 2916 498 2920 563
rect 2906 481 2908 483
rect 2925 481 2927 483
rect 2862 464 2864 476
rect 2881 474 2883 476
rect 2906 464 2908 476
rect 2862 462 2883 464
rect 2862 450 2864 453
rect 2881 450 2883 462
rect 2907 460 2908 464
rect 2925 463 2927 476
rect 2906 450 2908 460
rect 2926 459 2927 463
rect 2936 461 2942 463
rect 2925 450 2927 459
rect 2862 433 2864 445
rect 2881 437 2883 445
rect 2906 443 2908 445
rect 2925 437 2927 445
rect 2881 435 2927 437
rect 2940 433 2942 461
rect 2847 431 2942 433
rect 1343 427 1346 431
rect 1343 407 1346 423
rect 1354 419 1357 431
rect 2993 418 2997 563
rect 3052 514 3088 516
rect 3052 437 3054 514
rect 3067 485 3069 487
rect 3086 485 3088 514
rect 3113 502 3117 563
rect 3111 485 3113 487
rect 3130 485 3132 487
rect 3067 468 3069 480
rect 3086 478 3088 480
rect 3111 468 3113 480
rect 3130 468 3132 480
rect 3067 466 3088 468
rect 3067 454 3069 457
rect 3086 454 3088 466
rect 3112 464 3113 468
rect 3131 464 3132 468
rect 3141 465 3147 467
rect 3111 454 3113 464
rect 3130 454 3132 464
rect 3067 437 3069 449
rect 3086 441 3088 449
rect 3111 447 3113 449
rect 3130 441 3132 449
rect 3086 439 3132 441
rect 3145 437 3147 465
rect 3274 459 3278 563
rect 3235 447 3238 451
rect 3246 447 3249 451
rect 3052 435 3147 437
rect 3235 436 3238 440
rect 2993 417 3051 418
rect 1354 407 1357 415
rect 2892 413 3051 417
rect 1376 409 2339 413
rect 1343 395 1346 398
rect 1354 395 1357 398
rect 1376 382 1380 409
rect 1458 389 1462 409
rect 1570 392 1574 409
rect 1685 393 1689 409
rect 1807 394 1811 409
rect 1989 395 1993 409
rect 2101 397 2105 409
rect 2217 397 2221 409
rect 2335 398 2339 409
rect 2892 404 2896 413
rect 3047 404 3051 413
rect 2862 392 2865 396
rect 2873 392 2876 396
rect 2920 392 2923 395
rect 3017 392 3020 396
rect 3028 392 3031 396
rect 3075 392 3078 395
rect 1316 378 1380 382
rect 1429 379 1432 383
rect 1440 379 1443 383
rect 1487 379 1490 382
rect 1540 381 1543 385
rect 1551 381 1554 385
rect 1598 381 1601 384
rect 1656 381 1659 385
rect 1667 381 1670 385
rect 1714 381 1717 384
rect 1776 382 1779 386
rect 1787 382 1790 386
rect 1834 382 1837 385
rect 1958 383 1961 387
rect 1969 383 1972 387
rect 2016 383 2019 386
rect 2069 385 2072 389
rect 2080 385 2083 389
rect 2127 385 2130 388
rect 2185 385 2188 389
rect 2196 385 2199 389
rect 2243 385 2246 388
rect 2305 386 2308 390
rect 2316 386 2319 390
rect 2363 386 2366 389
rect 1316 356 1320 378
rect 1322 344 1325 348
rect 1333 344 1336 348
rect 1322 333 1325 337
rect 1322 313 1325 329
rect 1333 325 1336 337
rect 1333 313 1336 321
rect 1322 301 1325 304
rect 1333 301 1336 304
rect 1332 292 1333 295
rect 1328 280 1333 292
rect 1142 279 1364 280
rect 1144 275 1364 279
rect 981 270 1125 274
rect 981 263 985 270
rect 768 259 995 263
rect 991 247 995 259
rect 1121 258 1125 270
rect 1090 246 1093 250
rect 1101 246 1104 250
rect 1148 246 1151 249
rect 989 235 992 238
rect 1090 235 1093 239
rect 989 215 992 230
rect 1090 215 1093 231
rect 1101 227 1104 239
rect 1148 226 1151 241
rect 1101 215 1104 223
rect 989 196 992 211
rect 1148 207 1151 222
rect 1090 203 1093 206
rect 1101 203 1104 206
rect 1148 198 1151 202
rect 989 187 992 191
rect 987 175 991 176
rect 1124 175 1128 192
rect 1187 188 1191 275
rect 1187 184 1201 188
rect 1197 175 1201 184
rect 987 171 1201 175
rect 986 161 1122 165
rect 986 154 990 161
rect 768 150 997 154
rect 993 149 997 150
rect 990 138 993 141
rect 990 118 993 133
rect 990 99 993 114
rect 990 90 993 94
rect 1032 91 1036 161
rect 1118 158 1122 161
rect 1088 146 1091 150
rect 1099 146 1102 150
rect 1146 146 1149 149
rect 1088 135 1091 139
rect 1088 115 1091 131
rect 1099 127 1102 139
rect 1146 126 1149 141
rect 1099 115 1102 123
rect 1146 107 1149 122
rect 1088 103 1091 106
rect 1099 103 1102 106
rect 1146 98 1149 102
rect 1032 87 1123 91
rect 990 -8 993 79
rect 1119 69 1123 87
rect 1128 83 1132 95
rect 1197 83 1201 171
rect 1128 79 1201 83
rect 1089 57 1092 61
rect 1100 57 1103 61
rect 1147 57 1150 60
rect 1089 46 1092 50
rect 1089 26 1092 42
rect 1100 38 1103 50
rect 1147 37 1150 52
rect 1100 26 1103 34
rect 1147 18 1150 33
rect 1089 14 1092 17
rect 1100 14 1103 17
rect 1147 9 1150 13
rect 1124 -8 1128 5
rect 1197 -8 1201 79
rect 990 -11 1201 -8
rect 1124 -12 1201 -11
rect 1328 87 1333 275
rect 1376 211 1380 378
rect 1429 368 1432 372
rect 1429 348 1432 364
rect 1440 360 1443 372
rect 1487 359 1490 374
rect 1540 370 1543 374
rect 1440 348 1443 356
rect 1487 340 1490 355
rect 1540 350 1543 366
rect 1551 362 1554 374
rect 1598 361 1601 376
rect 1656 370 1659 374
rect 1551 350 1554 358
rect 1598 342 1601 357
rect 1656 350 1659 366
rect 1667 362 1670 374
rect 1714 361 1717 376
rect 1776 371 1779 375
rect 1667 350 1670 358
rect 1429 336 1432 339
rect 1440 336 1443 339
rect 1540 338 1543 341
rect 1551 338 1554 341
rect 1714 342 1717 357
rect 1776 351 1779 367
rect 1787 363 1790 375
rect 1834 362 1837 377
rect 1958 372 1961 376
rect 1787 351 1790 359
rect 1834 343 1837 358
rect 1958 352 1961 368
rect 1969 364 1972 376
rect 2016 363 2019 378
rect 2069 374 2072 378
rect 1969 352 1972 360
rect 2016 344 2019 359
rect 2069 354 2072 370
rect 2080 366 2083 378
rect 2127 365 2130 380
rect 2185 374 2188 378
rect 2080 354 2083 362
rect 2127 346 2130 361
rect 2185 354 2188 370
rect 2196 366 2199 378
rect 2243 365 2246 380
rect 2862 381 2865 385
rect 2305 375 2308 379
rect 2196 354 2199 362
rect 1656 338 1659 341
rect 1667 338 1670 341
rect 1776 339 1779 342
rect 1787 339 1790 342
rect 1958 340 1961 343
rect 1969 340 1972 343
rect 2069 342 2072 345
rect 2080 342 2083 345
rect 2243 346 2246 361
rect 2305 355 2308 371
rect 2316 367 2319 379
rect 2363 366 2366 381
rect 2316 355 2319 363
rect 2363 347 2366 362
rect 2862 361 2865 377
rect 2873 373 2876 385
rect 2920 372 2923 387
rect 3017 381 3020 385
rect 2873 361 2876 369
rect 2920 353 2923 368
rect 3017 361 3020 377
rect 3028 373 3031 385
rect 3075 372 3078 387
rect 3028 361 3031 369
rect 2862 349 2865 352
rect 2873 349 2876 352
rect 3075 353 3078 368
rect 3017 349 3020 352
rect 3028 349 3031 352
rect 2185 342 2188 345
rect 2196 342 2199 345
rect 2305 343 2308 346
rect 2316 343 2319 346
rect 2920 344 2923 348
rect 3075 344 3078 348
rect 3103 345 3107 419
rect 3235 416 3238 432
rect 3246 428 3249 440
rect 3246 416 3249 424
rect 3235 404 3238 407
rect 3246 404 3249 407
rect 3274 386 3278 455
rect 3587 526 3623 528
rect 3313 446 3316 450
rect 3324 446 3327 450
rect 3587 449 3589 526
rect 3602 497 3604 499
rect 3621 497 3623 526
rect 3651 513 3655 586
rect 3646 497 3648 499
rect 3665 497 3667 499
rect 3602 480 3604 492
rect 3621 490 3623 492
rect 3646 480 3648 492
rect 3602 478 3623 480
rect 3602 466 3604 469
rect 3621 466 3623 478
rect 3647 476 3648 480
rect 3665 479 3667 492
rect 3646 466 3648 476
rect 3666 475 3667 479
rect 3676 477 3682 479
rect 3665 466 3667 475
rect 3602 449 3604 461
rect 3621 453 3623 461
rect 3646 459 3648 461
rect 3665 453 3667 461
rect 3621 451 3667 453
rect 3680 449 3682 477
rect 3587 447 3682 449
rect 3313 435 3316 439
rect 3313 415 3316 431
rect 3324 427 3327 439
rect 3734 434 3738 586
rect 3856 585 4024 586
rect 3792 530 3828 532
rect 3792 453 3794 530
rect 3807 501 3809 503
rect 3826 501 3828 530
rect 3856 518 3860 585
rect 3851 501 3853 503
rect 3870 501 3872 503
rect 3807 484 3809 496
rect 3826 494 3828 496
rect 3851 484 3853 496
rect 3870 484 3872 496
rect 3807 482 3828 484
rect 3807 470 3809 473
rect 3826 470 3828 482
rect 3852 480 3853 484
rect 3871 480 3872 484
rect 3881 481 3887 483
rect 3851 470 3853 480
rect 3870 470 3872 480
rect 3807 453 3809 465
rect 3826 457 3828 465
rect 3851 463 3853 465
rect 3870 457 3872 465
rect 3826 455 3872 457
rect 3885 453 3887 481
rect 4020 475 4024 585
rect 4609 576 4613 722
rect 5233 717 5237 986
rect 5233 713 5294 717
rect 5172 697 5208 699
rect 5172 620 5174 697
rect 5187 668 5189 670
rect 5206 668 5208 697
rect 5233 685 5237 713
rect 5231 668 5233 670
rect 5250 668 5252 670
rect 5187 651 5189 663
rect 5206 661 5208 663
rect 5231 651 5233 663
rect 5250 651 5252 663
rect 5187 649 5208 651
rect 5187 637 5189 640
rect 5206 637 5208 649
rect 5232 647 5233 651
rect 5251 647 5252 651
rect 5261 648 5267 650
rect 5231 637 5233 647
rect 5250 637 5252 647
rect 5187 620 5189 632
rect 5206 624 5208 632
rect 5231 630 5233 632
rect 5250 624 5252 632
rect 5206 622 5252 624
rect 5265 620 5267 648
rect 5172 618 5267 620
rect 4609 575 4794 576
rect 4428 571 4794 575
rect 3975 463 3978 467
rect 3986 463 3989 467
rect 3792 451 3887 453
rect 3975 452 3978 456
rect 3324 415 3327 423
rect 3629 430 3791 434
rect 3629 420 3633 430
rect 3787 420 3791 430
rect 3602 408 3605 412
rect 3613 408 3616 412
rect 3660 408 3663 411
rect 3757 408 3760 412
rect 3768 408 3771 412
rect 3815 408 3818 411
rect 3313 403 3316 406
rect 3324 403 3327 406
rect 3602 397 3605 401
rect 3274 382 3298 386
rect 3294 367 3298 382
rect 3602 377 3605 393
rect 3613 389 3616 401
rect 3660 388 3663 403
rect 3757 397 3760 401
rect 3613 377 3616 385
rect 3660 369 3663 384
rect 3757 377 3760 393
rect 3768 389 3771 401
rect 3815 388 3818 403
rect 3768 377 3771 385
rect 3602 365 3605 368
rect 3613 365 3616 368
rect 3815 369 3818 384
rect 3757 365 3760 368
rect 3768 365 3771 368
rect 3660 360 3663 364
rect 3815 360 3818 364
rect 3292 352 3295 356
rect 3303 352 3306 356
rect 3635 347 3639 358
rect 3791 347 3795 354
rect 3849 347 3853 440
rect 3975 432 3978 448
rect 3986 444 3989 456
rect 3986 432 3989 440
rect 3975 420 3978 423
rect 3986 420 3989 423
rect 3970 347 3974 413
rect 4020 398 4024 471
rect 4366 537 4402 539
rect 4053 462 4056 466
rect 4064 462 4067 466
rect 4366 460 4368 537
rect 4381 508 4383 510
rect 4400 508 4402 537
rect 4428 525 4432 571
rect 4425 508 4427 510
rect 4444 508 4446 510
rect 4381 491 4383 503
rect 4400 501 4402 503
rect 4425 491 4427 503
rect 4381 489 4402 491
rect 4381 477 4383 480
rect 4400 477 4402 489
rect 4426 487 4427 491
rect 4444 490 4446 503
rect 4425 477 4427 487
rect 4445 486 4446 490
rect 4455 488 4461 490
rect 4444 477 4446 486
rect 4381 460 4383 472
rect 4400 464 4402 472
rect 4425 470 4427 472
rect 4444 464 4446 472
rect 4400 462 4446 464
rect 4459 460 4461 488
rect 4366 458 4461 460
rect 4053 451 4056 455
rect 4053 431 4056 447
rect 4064 443 4067 455
rect 4527 446 4531 571
rect 4571 541 4607 543
rect 4571 464 4573 541
rect 4586 512 4588 514
rect 4605 512 4607 541
rect 4633 529 4637 571
rect 4630 512 4632 514
rect 4649 512 4651 514
rect 4586 495 4588 507
rect 4605 505 4607 507
rect 4630 495 4632 507
rect 4649 495 4651 507
rect 4586 493 4607 495
rect 4586 481 4588 484
rect 4605 481 4607 493
rect 4631 491 4632 495
rect 4650 491 4651 495
rect 4660 492 4666 494
rect 4630 481 4632 491
rect 4649 481 4651 491
rect 4586 464 4588 476
rect 4605 468 4607 476
rect 4630 474 4632 476
rect 4649 468 4651 476
rect 4605 466 4651 468
rect 4664 464 4666 492
rect 4789 486 4794 571
rect 5290 568 5294 713
rect 5110 567 5294 568
rect 5311 567 5474 568
rect 5110 564 5474 567
rect 5110 563 5315 564
rect 4754 474 4757 478
rect 4765 474 4768 478
rect 4571 462 4666 464
rect 4754 463 4757 467
rect 4527 445 4570 446
rect 4064 431 4067 439
rect 4409 441 4570 445
rect 4409 431 4413 441
rect 4566 431 4570 441
rect 4053 419 4056 422
rect 4064 419 4067 422
rect 4381 419 4384 423
rect 4392 419 4395 423
rect 4439 419 4442 422
rect 4536 419 4539 423
rect 4547 419 4550 423
rect 4594 419 4597 422
rect 4381 408 4384 412
rect 4020 394 4042 398
rect 4038 383 4042 394
rect 4381 388 4384 404
rect 4392 400 4395 412
rect 4439 399 4442 414
rect 4536 408 4539 412
rect 4392 388 4395 396
rect 4439 380 4442 395
rect 4536 388 4539 404
rect 4547 400 4550 412
rect 4594 399 4597 414
rect 4547 388 4550 396
rect 4381 376 4384 379
rect 4392 376 4395 379
rect 4594 380 4597 395
rect 4536 376 4539 379
rect 4547 376 4550 379
rect 4032 368 4035 372
rect 4043 368 4046 372
rect 4439 371 4442 375
rect 4594 371 4597 375
rect 4411 361 4415 369
rect 4565 361 4569 365
rect 4032 357 4035 361
rect 1487 331 1490 335
rect 1598 333 1601 337
rect 1714 333 1717 337
rect 1834 334 1837 338
rect 2016 335 2019 339
rect 2127 337 2130 341
rect 2243 337 2246 341
rect 2363 338 2366 342
rect 1461 317 1465 327
rect 1572 317 1576 329
rect 1686 317 1690 329
rect 1808 317 1812 330
rect 1990 329 1994 331
rect 2101 329 2105 333
rect 2217 329 2221 333
rect 2337 329 2341 334
rect 2888 329 2892 342
rect 3046 329 3051 339
rect 3103 341 3227 345
rect 3292 341 3295 345
rect 3103 329 3107 341
rect 1873 324 3107 329
rect 1873 317 1878 324
rect 1403 312 1878 317
rect 1403 280 1408 312
rect 3180 293 3184 341
rect 3292 321 3295 337
rect 3303 333 3306 345
rect 3303 321 3306 329
rect 3569 343 3974 347
rect 3292 309 3295 312
rect 3303 309 3306 312
rect 3569 293 3573 343
rect 3970 325 3974 343
rect 4032 337 4035 353
rect 4043 349 4046 361
rect 4411 357 4569 361
rect 4043 337 4046 345
rect 4434 336 4437 357
rect 4627 336 4631 449
rect 4754 443 4757 459
rect 4765 455 4768 467
rect 4765 443 4768 451
rect 4754 431 4757 434
rect 4765 431 4768 434
rect 4750 336 4754 424
rect 4789 420 4794 482
rect 5046 531 5082 533
rect 4832 473 4835 477
rect 4843 473 4846 477
rect 4832 462 4835 466
rect 4832 442 4835 458
rect 4843 454 4846 466
rect 5046 454 5048 531
rect 5061 502 5063 504
rect 5080 502 5082 531
rect 5110 519 5114 563
rect 5105 502 5107 504
rect 5124 502 5126 504
rect 5061 485 5063 497
rect 5080 495 5082 497
rect 5105 485 5107 497
rect 5061 483 5082 485
rect 5061 471 5063 474
rect 5080 471 5082 483
rect 5106 481 5107 485
rect 5124 484 5126 497
rect 5105 471 5107 481
rect 5125 480 5126 484
rect 5135 482 5141 484
rect 5124 471 5126 480
rect 5061 454 5063 466
rect 5080 458 5082 466
rect 5105 464 5107 466
rect 5124 458 5126 466
rect 5080 456 5126 458
rect 5139 454 5141 482
rect 5046 452 5141 454
rect 4843 442 4846 450
rect 5157 445 5167 450
rect 5200 434 5205 563
rect 5251 535 5287 537
rect 5251 458 5253 535
rect 5266 506 5268 508
rect 5285 506 5287 535
rect 5311 523 5315 563
rect 5310 506 5312 508
rect 5329 506 5331 508
rect 5266 489 5268 501
rect 5285 499 5287 501
rect 5310 489 5312 501
rect 5329 489 5331 501
rect 5266 487 5287 489
rect 5266 475 5268 478
rect 5285 475 5287 487
rect 5311 485 5312 489
rect 5330 485 5331 489
rect 5340 486 5346 488
rect 5310 475 5312 485
rect 5329 475 5331 485
rect 5266 458 5268 470
rect 5285 462 5287 470
rect 5310 468 5312 470
rect 5329 462 5331 470
rect 5285 460 5331 462
rect 5344 458 5346 486
rect 5470 480 5474 564
rect 5434 468 5437 472
rect 5445 468 5448 472
rect 5251 456 5346 458
rect 5434 457 5437 461
rect 4832 430 4835 433
rect 4843 430 4846 433
rect 5089 429 5253 434
rect 5089 425 5094 429
rect 5248 425 5253 429
rect 4789 415 4819 420
rect 4814 394 4819 415
rect 5061 413 5064 417
rect 5072 413 5075 417
rect 5119 413 5122 416
rect 5216 413 5219 417
rect 5227 413 5230 417
rect 5274 413 5277 416
rect 5061 402 5064 406
rect 4811 379 4814 383
rect 4822 379 4825 383
rect 5061 382 5064 398
rect 5072 394 5075 406
rect 5119 393 5122 408
rect 5216 402 5219 406
rect 5072 382 5075 390
rect 5119 374 5122 389
rect 5216 382 5219 398
rect 5227 394 5230 406
rect 5274 393 5277 408
rect 5227 382 5230 390
rect 4811 368 4814 372
rect 4811 348 4814 364
rect 4822 360 4825 372
rect 5061 370 5064 373
rect 5072 370 5075 373
rect 5274 374 5277 389
rect 5216 370 5219 373
rect 5227 370 5230 373
rect 4822 348 4825 356
rect 5119 365 5122 369
rect 5094 352 5098 363
rect 5274 365 5277 369
rect 5245 352 5249 362
rect 5308 352 5312 443
rect 5434 437 5437 453
rect 5445 449 5448 461
rect 5445 437 5448 445
rect 5434 425 5437 428
rect 5445 425 5448 428
rect 5435 352 5439 417
rect 5470 411 5474 476
rect 5512 467 5515 471
rect 5523 467 5526 471
rect 5512 456 5515 460
rect 5512 436 5515 452
rect 5523 448 5526 460
rect 5523 436 5526 444
rect 5512 424 5515 427
rect 5523 424 5526 427
rect 5470 407 5497 411
rect 5493 388 5497 407
rect 5491 373 5494 377
rect 5502 373 5505 377
rect 5491 362 5494 366
rect 5065 348 5439 352
rect 4811 336 4814 339
rect 4822 336 4825 339
rect 4392 332 4754 336
rect 4032 325 4035 328
rect 4043 325 4046 328
rect 3970 321 4024 325
rect 3970 310 3974 321
rect 4392 310 4396 332
rect 4750 329 4754 332
rect 4750 327 4818 329
rect 4750 325 4822 327
rect 4750 318 4754 325
rect 5065 318 5069 348
rect 4750 314 5069 318
rect 5435 320 5439 348
rect 5491 342 5494 358
rect 5502 354 5505 366
rect 5502 342 5505 350
rect 5491 330 5494 333
rect 5502 330 5505 333
rect 5501 320 5505 322
rect 5435 316 5505 320
rect 3970 306 4396 310
rect 3180 289 3573 293
rect 1395 275 1408 280
rect 1376 207 2343 211
rect 1328 82 1362 87
rect 1124 -45 1128 -12
rect 1328 -64 1333 82
rect 1376 30 1380 207
rect 1461 189 1465 207
rect 1572 191 1576 207
rect 1688 191 1692 207
rect 1808 192 1812 207
rect 1991 193 1995 207
rect 2104 195 2108 207
rect 2219 195 2223 207
rect 2339 196 2343 207
rect 1432 177 1435 181
rect 1443 177 1446 181
rect 1490 177 1493 180
rect 1543 179 1546 183
rect 1554 179 1557 183
rect 1601 179 1604 182
rect 1659 179 1662 183
rect 1670 179 1673 183
rect 1717 179 1720 182
rect 1779 180 1782 184
rect 1790 180 1793 184
rect 1837 180 1840 183
rect 1961 181 1964 185
rect 1972 181 1975 185
rect 2019 181 2022 184
rect 2072 183 2075 187
rect 2083 183 2086 187
rect 2130 183 2133 186
rect 2188 183 2191 187
rect 2199 183 2202 187
rect 2246 183 2249 186
rect 2308 184 2311 188
rect 2319 184 2322 188
rect 2366 184 2369 187
rect 1432 166 1435 170
rect 1432 146 1435 162
rect 1443 158 1446 170
rect 1490 157 1493 172
rect 1543 168 1546 172
rect 1443 146 1446 154
rect 1490 138 1493 153
rect 1543 148 1546 164
rect 1554 160 1557 172
rect 1601 159 1604 174
rect 1659 168 1662 172
rect 1554 148 1557 156
rect 1601 140 1604 155
rect 1659 148 1662 164
rect 1670 160 1673 172
rect 1717 159 1720 174
rect 1779 169 1782 173
rect 1670 148 1673 156
rect 1432 134 1435 137
rect 1443 134 1446 137
rect 1543 136 1546 139
rect 1554 136 1557 139
rect 1717 140 1720 155
rect 1779 149 1782 165
rect 1790 161 1793 173
rect 1837 160 1840 175
rect 1961 170 1964 174
rect 1790 149 1793 157
rect 1837 141 1840 156
rect 1961 150 1964 166
rect 1972 162 1975 174
rect 2019 161 2022 176
rect 2072 172 2075 176
rect 1972 150 1975 158
rect 2019 142 2022 157
rect 2072 152 2075 168
rect 2083 164 2086 176
rect 2130 163 2133 178
rect 2188 172 2191 176
rect 2083 152 2086 160
rect 2130 144 2133 159
rect 2188 152 2191 168
rect 2199 164 2202 176
rect 2246 163 2249 178
rect 2308 173 2311 177
rect 2199 152 2202 160
rect 1659 136 1662 139
rect 1670 136 1673 139
rect 1779 137 1782 140
rect 1790 137 1793 140
rect 1961 138 1964 141
rect 1972 138 1975 141
rect 2072 140 2075 143
rect 2083 140 2086 143
rect 2246 144 2249 159
rect 2308 153 2311 169
rect 2319 165 2322 177
rect 2366 164 2369 179
rect 2319 153 2322 161
rect 2366 145 2369 160
rect 2188 140 2191 143
rect 2199 140 2202 143
rect 2308 141 2311 144
rect 2319 141 2322 144
rect 1490 129 1493 133
rect 1601 131 1604 135
rect 1717 131 1720 135
rect 1837 132 1840 136
rect 2019 133 2022 137
rect 2130 135 2133 139
rect 2246 135 2249 139
rect 2366 136 2369 140
rect 1464 120 1468 125
rect 1574 120 1578 127
rect 1691 120 1695 127
rect 1811 120 1815 128
rect 1993 120 1997 129
rect 2105 120 2109 131
rect 2220 120 2224 131
rect 2341 120 2345 132
rect 1401 115 2345 120
rect 1401 87 1406 115
rect 1393 82 1406 87
rect 3558 47 4112 51
rect 3558 30 3562 47
rect 1376 26 3562 30
rect 3631 28 3635 47
rect 1328 -69 1362 -64
rect 1328 -205 1333 -69
rect 1376 -119 1380 26
rect 1486 12 1490 26
rect 1597 14 1601 26
rect 1712 14 1716 26
rect 1834 15 1838 26
rect 2016 16 2020 26
rect 2128 18 2132 26
rect 2245 18 2249 26
rect 2364 19 2368 26
rect 1457 1 1460 4
rect 1468 1 1471 4
rect 1515 1 1518 3
rect 1568 1 1571 6
rect 1457 -11 1460 -5
rect 1457 -31 1460 -15
rect 1468 -19 1471 -5
rect 1515 -20 1518 -3
rect 1579 1 1582 6
rect 1626 1 1629 5
rect 1684 1 1687 6
rect 1695 1 1698 6
rect 1742 0 1745 2
rect 1568 -9 1571 -5
rect 1468 -31 1471 -23
rect 1515 -39 1518 -24
rect 1568 -29 1571 -13
rect 1579 -17 1582 -5
rect 1626 -18 1629 -3
rect 1684 -9 1687 -2
rect 1579 -29 1582 -21
rect 1626 -37 1629 -22
rect 1684 -29 1687 -13
rect 1695 -17 1698 -2
rect 1804 2 1807 7
rect 1815 2 1818 7
rect 1862 0 1865 6
rect 1986 4 1989 8
rect 1997 4 2000 8
rect 2044 4 2047 7
rect 1742 -18 1745 -4
rect 1804 -8 1807 -1
rect 1695 -29 1698 -21
rect 1457 -43 1460 -40
rect 1468 -43 1471 -40
rect 1568 -41 1571 -38
rect 1579 -41 1582 -38
rect 1742 -37 1745 -22
rect 1804 -28 1807 -12
rect 1815 -16 1818 -1
rect 1862 -17 1865 -4
rect 1986 -7 1989 1
rect 1815 -28 1818 -20
rect 1862 -36 1865 -21
rect 1986 -27 1989 -11
rect 1997 -15 2000 1
rect 2097 6 2100 10
rect 2108 6 2111 10
rect 2155 6 2158 9
rect 2213 6 2216 10
rect 2224 6 2227 10
rect 2271 6 2274 9
rect 2333 7 2336 11
rect 2344 7 2347 11
rect 2391 7 2394 10
rect 2044 -16 2047 0
rect 2097 -5 2100 3
rect 1997 -27 2000 -19
rect 2044 -35 2047 -20
rect 2097 -25 2100 -9
rect 2108 -13 2111 3
rect 2155 -14 2158 3
rect 2213 -5 2216 3
rect 2108 -25 2111 -17
rect 2155 -33 2158 -18
rect 2213 -25 2216 -9
rect 2224 -13 2227 3
rect 2271 -14 2274 3
rect 2333 -4 2336 3
rect 2224 -25 2227 -17
rect 1684 -41 1687 -38
rect 1695 -41 1698 -38
rect 1804 -40 1807 -37
rect 1815 -40 1818 -37
rect 1986 -39 1989 -36
rect 1997 -39 2000 -36
rect 2097 -37 2100 -34
rect 2108 -37 2111 -34
rect 2271 -33 2274 -18
rect 2333 -24 2336 -8
rect 2344 -12 2347 3
rect 2391 -13 2394 3
rect 2344 -24 2347 -16
rect 2391 -32 2394 -17
rect 2213 -37 2216 -34
rect 2224 -37 2227 -34
rect 2333 -36 2336 -33
rect 2344 -36 2347 -33
rect 1515 -48 1518 -44
rect 1626 -46 1629 -42
rect 1742 -46 1745 -42
rect 1862 -45 1865 -41
rect 2044 -44 2047 -40
rect 2155 -42 2158 -38
rect 2271 -42 2274 -38
rect 2391 -41 2394 -37
rect 1489 -55 1493 -52
rect 1600 -55 1604 -50
rect 1715 -55 1719 -50
rect 1836 -55 1840 -49
rect 2018 -55 2022 -48
rect 2129 -55 2133 -46
rect 2245 -55 2249 -46
rect 2366 -55 2370 -45
rect 1401 -60 2370 -55
rect 1401 -64 1406 -60
rect 1393 -69 1406 -64
rect 1376 -123 2128 -119
rect 1755 -129 1759 -123
rect 1871 -130 1875 -123
rect 2004 -131 2009 -123
rect 2124 -131 2128 -123
rect 1724 -141 1727 -137
rect 1735 -141 1738 -137
rect 1782 -141 1785 -138
rect 1842 -142 1845 -138
rect 1853 -142 1856 -138
rect 1900 -142 1903 -139
rect 1975 -142 1978 -138
rect 1986 -142 1989 -138
rect 2033 -142 2036 -139
rect 1724 -152 1727 -148
rect 1724 -172 1727 -156
rect 1735 -160 1738 -148
rect 1782 -161 1785 -146
rect 1842 -153 1845 -149
rect 1735 -172 1738 -164
rect 1782 -180 1785 -165
rect 1842 -173 1845 -157
rect 1853 -161 1856 -149
rect 1900 -162 1903 -147
rect 2094 -143 2097 -139
rect 2105 -143 2108 -139
rect 2152 -143 2155 -140
rect 1975 -153 1978 -149
rect 1853 -173 1856 -165
rect 1724 -184 1727 -181
rect 1735 -184 1738 -181
rect 1900 -181 1903 -166
rect 1975 -173 1978 -157
rect 1986 -161 1989 -149
rect 2033 -162 2036 -147
rect 2094 -154 2097 -150
rect 1986 -173 1989 -165
rect 1842 -185 1845 -182
rect 1853 -185 1856 -182
rect 1782 -189 1785 -185
rect 2033 -181 2036 -166
rect 2094 -174 2097 -158
rect 2105 -162 2108 -150
rect 2152 -163 2155 -148
rect 2105 -174 2108 -166
rect 1975 -185 1978 -182
rect 1986 -185 1989 -182
rect 2152 -182 2155 -167
rect 2094 -186 2097 -183
rect 2105 -186 2108 -183
rect 1900 -190 1903 -186
rect 2033 -190 2036 -186
rect 2152 -191 2155 -187
rect 1754 -205 1758 -192
rect 1873 -205 1877 -196
rect 2006 -205 2010 -195
rect 2122 -205 2126 -195
rect 1328 -210 2281 -205
rect 2276 -211 2281 -210
rect 2276 -215 2782 -211
rect 2773 -598 2777 -215
rect 2818 -574 2822 26
rect 3537 -195 3541 26
rect 3592 16 3595 20
rect 3603 16 3606 20
rect 3592 5 3595 9
rect 3592 -15 3595 1
rect 3603 -3 3606 9
rect 3603 -15 3606 -7
rect 3592 -27 3595 -24
rect 3603 -27 3606 -24
rect 3596 -145 3600 -33
rect 3631 -54 3635 24
rect 3670 15 3673 19
rect 3681 15 3684 19
rect 3670 4 3673 8
rect 3670 -16 3673 0
rect 3681 -4 3684 8
rect 3681 -16 3684 -8
rect 3670 -28 3673 -25
rect 3681 -28 3684 -25
rect 3631 -57 3658 -54
rect 3654 -64 3658 -57
rect 3649 -79 3652 -75
rect 3660 -79 3663 -75
rect 3649 -90 3652 -86
rect 3649 -110 3652 -94
rect 3660 -98 3663 -86
rect 3660 -110 3663 -102
rect 3649 -122 3652 -119
rect 3660 -122 3663 -119
rect 3656 -145 3660 -131
rect 3596 -149 3660 -145
rect 3656 -176 3660 -149
rect 3681 -176 3685 -35
rect 3839 -99 3843 47
rect 3810 -111 3813 -107
rect 3821 -111 3824 -107
rect 3810 -122 3813 -118
rect 3810 -142 3813 -126
rect 3821 -130 3824 -118
rect 3839 -122 3843 -103
rect 3888 -112 3891 -108
rect 3899 -112 3902 -108
rect 3839 -126 3850 -122
rect 3888 -123 3891 -119
rect 3821 -142 3824 -134
rect 3810 -154 3813 -151
rect 3821 -154 3824 -151
rect 3815 -176 3819 -162
rect 3656 -180 3819 -176
rect 3537 -199 3653 -195
rect 2831 -215 3484 -211
rect 3480 -411 3484 -215
rect 3649 -248 3653 -199
rect 3605 -260 3608 -256
rect 3616 -260 3619 -256
rect 3605 -271 3608 -267
rect 3605 -291 3608 -275
rect 3616 -279 3619 -267
rect 3616 -291 3619 -283
rect 3605 -303 3608 -300
rect 3616 -303 3619 -300
rect 3610 -411 3614 -311
rect 3649 -336 3653 -252
rect 3683 -261 3686 -257
rect 3694 -261 3697 -257
rect 3683 -272 3686 -268
rect 3683 -292 3686 -276
rect 3694 -280 3697 -268
rect 3815 -270 3819 -180
rect 3846 -179 3850 -126
rect 3888 -143 3891 -127
rect 3899 -131 3902 -119
rect 3899 -143 3902 -135
rect 4108 -136 4112 47
rect 4104 -148 4107 -145
rect 3888 -155 3891 -152
rect 3899 -155 3902 -152
rect 3846 -183 3875 -179
rect 3871 -191 3875 -183
rect 3867 -206 3870 -202
rect 3878 -206 3881 -202
rect 3867 -217 3870 -213
rect 3867 -237 3870 -221
rect 3878 -225 3881 -213
rect 3878 -237 3881 -229
rect 3867 -249 3870 -246
rect 3878 -249 3881 -246
rect 3874 -269 3878 -257
rect 3904 -269 3908 -162
rect 4104 -168 4107 -153
rect 4104 -187 4107 -172
rect 4104 -196 4107 -192
rect 3874 -270 3908 -269
rect 3815 -273 3908 -270
rect 3815 -274 3878 -273
rect 3694 -292 3697 -284
rect 3683 -304 3686 -301
rect 3694 -304 3697 -301
rect 3649 -340 3670 -336
rect 3662 -355 3665 -351
rect 3673 -355 3676 -351
rect 3662 -366 3665 -362
rect 3662 -386 3665 -370
rect 3673 -374 3676 -362
rect 3673 -386 3676 -378
rect 3662 -398 3665 -395
rect 3673 -398 3676 -395
rect 3669 -411 3673 -406
rect 3694 -411 3698 -311
rect 3874 -411 3878 -274
rect 4106 -411 4110 -207
rect 3480 -415 4110 -411
rect 2818 -578 3643 -574
rect 2841 -580 2845 -578
rect 2837 -592 2840 -589
rect 2773 -602 2801 -598
rect 2797 -643 2801 -602
rect 2837 -612 2840 -597
rect 2837 -631 2840 -616
rect 2837 -640 2840 -636
rect 2797 -649 2821 -643
rect 2864 -823 2868 -578
rect 2911 -699 2915 -578
rect 3004 -580 3008 -578
rect 3002 -592 3005 -589
rect 3002 -612 3005 -597
rect 3002 -631 3005 -616
rect 3002 -640 3005 -636
rect 3085 -694 3089 -578
rect 3183 -579 3187 -578
rect 3179 -591 3182 -588
rect 3179 -611 3182 -596
rect 3179 -630 3182 -615
rect 3179 -639 3182 -635
rect 3275 -698 3279 -578
rect 3358 -580 3362 -578
rect 3354 -592 3357 -589
rect 3354 -612 3357 -597
rect 3354 -631 3357 -616
rect 3354 -640 3357 -636
rect 3457 -694 3461 -578
rect 3639 -604 3643 -578
rect 4198 -581 4638 -577
rect 4198 -604 4202 -581
rect 3639 -608 4202 -604
rect 3754 -625 3758 -608
rect 3752 -637 3755 -634
rect 3752 -657 3755 -642
rect 3752 -676 3755 -661
rect 3752 -685 3755 -681
rect 3053 -706 3056 -702
rect 3064 -706 3067 -702
rect 3111 -706 3114 -703
rect 3427 -706 3430 -702
rect 3438 -706 3441 -702
rect 3485 -706 3488 -703
rect 2882 -711 2885 -707
rect 2893 -711 2896 -707
rect 2940 -711 2943 -708
rect 3246 -710 3249 -706
rect 3257 -710 3260 -706
rect 3304 -710 3307 -707
rect 2882 -722 2885 -718
rect 2882 -742 2885 -726
rect 2893 -730 2896 -718
rect 2940 -731 2943 -716
rect 3053 -717 3056 -713
rect 2893 -742 2896 -734
rect 2940 -750 2943 -735
rect 3053 -737 3056 -721
rect 3064 -725 3067 -713
rect 3111 -726 3114 -711
rect 3246 -721 3249 -717
rect 3064 -737 3067 -729
rect 3111 -745 3114 -730
rect 3246 -741 3249 -725
rect 3257 -729 3260 -717
rect 3304 -730 3307 -715
rect 3427 -717 3430 -713
rect 3257 -741 3260 -733
rect 3053 -749 3056 -746
rect 3064 -749 3067 -746
rect 3304 -749 3307 -734
rect 3427 -737 3430 -721
rect 3438 -725 3441 -713
rect 3485 -726 3488 -711
rect 3438 -737 3441 -729
rect 3485 -745 3488 -730
rect 3427 -749 3430 -746
rect 3438 -749 3441 -746
rect 2882 -754 2885 -751
rect 2893 -754 2896 -751
rect 3111 -754 3114 -750
rect 3246 -753 3249 -750
rect 3257 -753 3260 -750
rect 3485 -754 3488 -750
rect 2940 -759 2943 -755
rect 3304 -758 3307 -754
rect 2913 -771 2917 -764
rect 3085 -771 3089 -759
rect 3277 -771 3281 -763
rect 3458 -770 3462 -759
rect 3737 -770 3741 -696
rect 3458 -771 3741 -770
rect 2913 -774 3741 -771
rect 2864 -827 3049 -823
rect 2864 -1016 2868 -827
rect 3045 -838 3049 -827
rect 3014 -850 3017 -846
rect 3025 -850 3028 -846
rect 3072 -850 3075 -847
rect 3014 -861 3017 -857
rect 3014 -881 3017 -865
rect 3025 -869 3028 -857
rect 3072 -870 3075 -855
rect 3025 -881 3028 -873
rect 3072 -889 3075 -874
rect 3014 -893 3017 -890
rect 3025 -893 3028 -890
rect 3072 -898 3075 -894
rect 3047 -909 3051 -902
rect 3113 -909 3116 -774
rect 3047 -912 3116 -909
rect 2864 -1020 3052 -1016
rect 2864 -1194 2868 -1020
rect 3048 -1036 3052 -1020
rect 3018 -1048 3021 -1044
rect 3029 -1048 3032 -1044
rect 3076 -1048 3079 -1045
rect 3018 -1059 3021 -1055
rect 3018 -1079 3021 -1063
rect 3029 -1067 3032 -1055
rect 3076 -1068 3079 -1053
rect 3029 -1079 3032 -1071
rect 3076 -1087 3079 -1072
rect 3018 -1091 3021 -1088
rect 3029 -1091 3032 -1088
rect 3076 -1096 3079 -1092
rect 3048 -1113 3052 -1100
rect 3113 -1113 3116 -912
rect 3793 -837 3797 -608
rect 3816 -621 3852 -619
rect 3816 -698 3818 -621
rect 3831 -650 3833 -648
rect 3850 -650 3852 -621
rect 3878 -633 3883 -608
rect 4003 -626 4007 -608
rect 4000 -638 4003 -635
rect 3875 -650 3877 -648
rect 3894 -650 3896 -648
rect 3831 -667 3833 -655
rect 3850 -657 3852 -655
rect 3875 -667 3877 -655
rect 3831 -669 3852 -667
rect 3831 -681 3833 -678
rect 3850 -681 3852 -669
rect 3876 -671 3877 -667
rect 3894 -668 3896 -655
rect 4000 -658 4003 -643
rect 3875 -681 3877 -671
rect 3895 -672 3896 -668
rect 3905 -670 3911 -668
rect 3894 -681 3896 -672
rect 3831 -698 3833 -686
rect 3850 -694 3852 -686
rect 3875 -688 3877 -686
rect 3894 -694 3896 -686
rect 3850 -696 3896 -694
rect 3909 -698 3911 -670
rect 4000 -677 4003 -662
rect 4000 -686 4003 -682
rect 3816 -700 3911 -698
rect 3793 -841 3899 -837
rect 3793 -1015 3797 -841
rect 3895 -870 3899 -841
rect 4006 -843 4010 -710
rect 4038 -751 4042 -608
rect 4064 -622 4100 -620
rect 4064 -699 4066 -622
rect 4079 -651 4081 -649
rect 4098 -651 4100 -622
rect 4125 -634 4129 -608
rect 4247 -617 4251 -581
rect 4307 -613 4343 -611
rect 4243 -629 4246 -626
rect 4243 -649 4246 -634
rect 4123 -651 4125 -649
rect 4142 -651 4144 -649
rect 4079 -668 4081 -656
rect 4098 -658 4100 -656
rect 4123 -668 4125 -656
rect 4142 -668 4144 -656
rect 4243 -668 4246 -653
rect 4079 -670 4100 -668
rect 4079 -682 4081 -679
rect 4098 -682 4100 -670
rect 4124 -672 4125 -668
rect 4143 -672 4144 -668
rect 4153 -671 4159 -669
rect 4123 -682 4125 -672
rect 4142 -682 4144 -672
rect 4079 -699 4081 -687
rect 4098 -695 4100 -687
rect 4123 -689 4125 -687
rect 4142 -695 4144 -687
rect 4098 -697 4144 -695
rect 4157 -699 4159 -671
rect 4243 -677 4246 -673
rect 4307 -690 4309 -613
rect 4322 -642 4324 -640
rect 4341 -642 4343 -613
rect 4363 -625 4367 -581
rect 4514 -612 4518 -581
rect 4576 -608 4612 -606
rect 4512 -624 4515 -621
rect 4366 -642 4368 -640
rect 4385 -642 4387 -640
rect 4512 -644 4515 -629
rect 4322 -659 4324 -647
rect 4341 -649 4343 -647
rect 4366 -659 4368 -647
rect 4385 -659 4387 -647
rect 4322 -661 4343 -659
rect 4322 -673 4324 -670
rect 4341 -673 4343 -661
rect 4367 -663 4368 -659
rect 4386 -663 4387 -659
rect 4396 -662 4402 -660
rect 4366 -673 4368 -663
rect 4385 -673 4387 -663
rect 4322 -690 4324 -678
rect 4341 -686 4343 -678
rect 4366 -680 4368 -678
rect 4385 -686 4387 -678
rect 4341 -688 4387 -686
rect 4400 -690 4402 -662
rect 4512 -663 4515 -648
rect 4512 -672 4515 -668
rect 4576 -685 4578 -608
rect 4591 -637 4593 -635
rect 4610 -637 4612 -608
rect 4634 -620 4638 -581
rect 4635 -637 4637 -635
rect 4654 -637 4656 -635
rect 4591 -654 4593 -642
rect 4610 -644 4612 -642
rect 4635 -654 4637 -642
rect 4654 -654 4656 -642
rect 4591 -656 4612 -654
rect 4591 -668 4593 -665
rect 4610 -668 4612 -656
rect 4636 -658 4637 -654
rect 4655 -658 4656 -654
rect 4665 -657 4671 -655
rect 4635 -668 4637 -658
rect 4654 -668 4656 -658
rect 4591 -685 4593 -673
rect 4610 -681 4612 -673
rect 4635 -675 4637 -673
rect 4654 -681 4656 -673
rect 4610 -683 4656 -681
rect 4669 -685 4671 -657
rect 4576 -687 4671 -685
rect 4307 -692 4402 -690
rect 4064 -701 4159 -699
rect 4038 -755 4493 -751
rect 4085 -767 4088 -763
rect 4096 -767 4099 -763
rect 4143 -767 4146 -764
rect 4085 -778 4088 -774
rect 4085 -798 4088 -782
rect 4096 -786 4099 -774
rect 4143 -787 4146 -772
rect 4335 -775 4339 -755
rect 4489 -767 4493 -755
rect 4461 -779 4464 -775
rect 4472 -779 4475 -775
rect 4519 -779 4522 -776
rect 4305 -787 4308 -783
rect 4316 -787 4319 -783
rect 4363 -787 4366 -784
rect 4096 -798 4099 -790
rect 4143 -806 4146 -791
rect 4461 -790 4464 -786
rect 4305 -798 4308 -794
rect 4085 -810 4088 -807
rect 4096 -810 4099 -807
rect 4143 -815 4146 -811
rect 4305 -818 4308 -802
rect 4316 -806 4319 -794
rect 4363 -807 4366 -792
rect 4316 -818 4319 -810
rect 4461 -810 4464 -794
rect 4472 -798 4475 -786
rect 4519 -799 4522 -784
rect 4472 -810 4475 -802
rect 4116 -843 4120 -819
rect 4363 -826 4366 -811
rect 4519 -818 4522 -803
rect 4461 -822 4464 -819
rect 4472 -822 4475 -819
rect 4305 -830 4308 -827
rect 4316 -830 4319 -827
rect 4519 -827 4522 -823
rect 4363 -835 4366 -831
rect 4336 -843 4340 -839
rect 4492 -843 4496 -831
rect 4006 -847 4496 -843
rect 3864 -882 3867 -878
rect 3875 -882 3878 -878
rect 3922 -882 3925 -879
rect 3864 -893 3867 -889
rect 3864 -913 3867 -897
rect 3875 -901 3878 -889
rect 3922 -902 3925 -887
rect 3875 -913 3878 -905
rect 3922 -921 3925 -906
rect 3864 -925 3867 -922
rect 3875 -925 3878 -922
rect 3922 -930 3925 -926
rect 3895 -940 3899 -935
rect 4006 -940 4010 -847
rect 3895 -944 4010 -940
rect 4006 -1004 4010 -944
rect 4844 -965 5264 -961
rect 3793 -1019 4238 -1015
rect 3905 -1056 3909 -1019
rect 3877 -1068 3880 -1064
rect 3888 -1068 3891 -1064
rect 3935 -1068 3938 -1065
rect 3877 -1079 3880 -1075
rect 3877 -1099 3880 -1083
rect 3888 -1087 3891 -1075
rect 3935 -1088 3938 -1073
rect 3888 -1099 3891 -1091
rect 3935 -1107 3938 -1092
rect 3877 -1111 3880 -1108
rect 3888 -1111 3891 -1108
rect 3048 -1116 3116 -1113
rect 3935 -1116 3938 -1112
rect 3095 -1187 3098 -1116
rect 3907 -1125 3911 -1120
rect 4006 -1125 4010 -1030
rect 4234 -1039 4238 -1019
rect 4205 -1051 4208 -1047
rect 4216 -1051 4219 -1047
rect 4263 -1051 4266 -1048
rect 4205 -1062 4208 -1058
rect 4205 -1082 4208 -1066
rect 4216 -1070 4219 -1058
rect 4263 -1071 4266 -1056
rect 4216 -1082 4219 -1074
rect 4263 -1090 4266 -1075
rect 4205 -1094 4208 -1091
rect 4216 -1094 4219 -1091
rect 4263 -1099 4266 -1095
rect 4242 -1125 4246 -1103
rect 3907 -1129 4246 -1125
rect 2864 -1198 3386 -1194
rect 2864 -1211 2868 -1198
rect 2862 -1223 2865 -1220
rect 2862 -1243 2865 -1228
rect 2862 -1262 2865 -1247
rect 2862 -1271 2865 -1267
rect 2913 -1319 2917 -1198
rect 3030 -1211 3034 -1198
rect 3207 -1210 3211 -1198
rect 3382 -1211 3386 -1198
rect 3027 -1223 3030 -1220
rect 3204 -1222 3207 -1219
rect 3379 -1223 3382 -1220
rect 3027 -1243 3030 -1228
rect 3204 -1242 3207 -1227
rect 3379 -1243 3382 -1228
rect 3027 -1262 3030 -1247
rect 3204 -1261 3207 -1246
rect 3379 -1262 3382 -1247
rect 3027 -1271 3030 -1267
rect 3204 -1270 3207 -1266
rect 3379 -1271 3382 -1267
rect 2913 -1323 3640 -1319
rect 2936 -1330 2940 -1323
rect 3107 -1325 3111 -1323
rect 3299 -1329 3303 -1323
rect 3482 -1325 3486 -1323
rect 3078 -1337 3081 -1333
rect 3089 -1337 3092 -1333
rect 3136 -1337 3139 -1334
rect 3452 -1337 3455 -1333
rect 3463 -1337 3466 -1333
rect 3510 -1337 3513 -1334
rect 2907 -1342 2910 -1338
rect 2918 -1342 2921 -1338
rect 2965 -1342 2968 -1339
rect 3271 -1341 3274 -1337
rect 3282 -1341 3285 -1337
rect 3329 -1341 3332 -1338
rect 2907 -1353 2910 -1349
rect 2907 -1373 2910 -1357
rect 2918 -1361 2921 -1349
rect 2965 -1362 2968 -1347
rect 3078 -1348 3081 -1344
rect 2918 -1373 2921 -1365
rect 2965 -1381 2968 -1366
rect 3078 -1368 3081 -1352
rect 3089 -1356 3092 -1344
rect 3136 -1357 3139 -1342
rect 3271 -1352 3274 -1348
rect 3089 -1368 3092 -1360
rect 3136 -1376 3139 -1361
rect 3271 -1372 3274 -1356
rect 3282 -1360 3285 -1348
rect 3329 -1361 3332 -1346
rect 3452 -1348 3455 -1344
rect 3282 -1372 3285 -1364
rect 3078 -1380 3081 -1377
rect 3089 -1380 3092 -1377
rect 3329 -1380 3332 -1365
rect 3452 -1368 3455 -1352
rect 3463 -1356 3466 -1344
rect 3510 -1357 3513 -1342
rect 3463 -1368 3466 -1360
rect 3510 -1376 3513 -1361
rect 3452 -1380 3455 -1377
rect 3463 -1380 3466 -1377
rect 2907 -1385 2910 -1382
rect 2918 -1385 2921 -1382
rect 3136 -1385 3139 -1381
rect 3271 -1384 3274 -1381
rect 3282 -1384 3285 -1381
rect 3510 -1385 3513 -1381
rect 2965 -1390 2968 -1386
rect 3329 -1389 3332 -1385
rect 2939 -1398 2943 -1395
rect 3110 -1398 3114 -1390
rect 3303 -1398 3307 -1394
rect 3484 -1398 3488 -1390
rect 2939 -1402 3488 -1398
rect 3484 -1944 3488 -1402
rect 3636 -1469 3640 -1323
rect 3636 -1473 4055 -1469
rect 3636 -1740 3640 -1473
rect 3705 -1526 3710 -1473
rect 3664 -1538 3667 -1534
rect 3675 -1538 3678 -1534
rect 3664 -1549 3667 -1545
rect 3664 -1569 3667 -1553
rect 3675 -1557 3678 -1545
rect 3675 -1569 3678 -1561
rect 3664 -1581 3667 -1578
rect 3675 -1581 3678 -1578
rect 3671 -1701 3675 -1590
rect 3705 -1617 3710 -1530
rect 3742 -1539 3745 -1535
rect 3753 -1539 3756 -1535
rect 3742 -1550 3745 -1546
rect 3742 -1570 3745 -1554
rect 3753 -1558 3756 -1546
rect 3753 -1570 3756 -1562
rect 4051 -1572 4055 -1473
rect 4844 -1572 4848 -965
rect 5045 -992 5049 -965
rect 5260 -993 5264 -965
rect 5015 -1004 5018 -1000
rect 5026 -1004 5029 -1000
rect 5073 -1004 5076 -1001
rect 5232 -1005 5235 -1001
rect 5243 -1005 5246 -1001
rect 5290 -1005 5293 -1002
rect 5015 -1015 5018 -1011
rect 5015 -1035 5018 -1019
rect 5026 -1023 5029 -1011
rect 5073 -1024 5076 -1009
rect 5232 -1016 5235 -1012
rect 5026 -1035 5029 -1027
rect 5073 -1043 5076 -1028
rect 5232 -1036 5235 -1020
rect 5243 -1024 5246 -1012
rect 5290 -1025 5293 -1010
rect 5243 -1036 5246 -1028
rect 5015 -1047 5018 -1044
rect 5026 -1047 5029 -1044
rect 5290 -1044 5293 -1029
rect 5232 -1048 5235 -1045
rect 5243 -1048 5246 -1045
rect 5073 -1052 5076 -1048
rect 5290 -1053 5293 -1049
rect 5046 -1065 5050 -1057
rect 5258 -1065 5262 -1058
rect 4051 -1576 4848 -1572
rect 5004 -1069 5262 -1065
rect 3742 -1582 3745 -1579
rect 3753 -1582 3756 -1579
rect 3705 -1621 3731 -1617
rect 3705 -1622 3726 -1621
rect 3721 -1633 3724 -1629
rect 3732 -1633 3735 -1629
rect 3721 -1644 3724 -1640
rect 3721 -1664 3724 -1648
rect 3732 -1652 3735 -1640
rect 3732 -1664 3735 -1656
rect 3721 -1676 3724 -1673
rect 3732 -1676 3735 -1673
rect 3729 -1701 3733 -1685
rect 3757 -1701 3761 -1589
rect 4051 -1636 4055 -1576
rect 4570 -1623 4574 -1576
rect 4566 -1635 4569 -1632
rect 4009 -1648 4012 -1644
rect 4020 -1648 4023 -1644
rect 4009 -1659 4012 -1655
rect 4009 -1679 4012 -1663
rect 4020 -1667 4023 -1655
rect 4020 -1679 4023 -1671
rect 4009 -1691 4012 -1688
rect 4020 -1691 4023 -1688
rect 3671 -1705 3908 -1701
rect 3636 -1744 3714 -1740
rect 3710 -1770 3714 -1744
rect 3674 -1782 3677 -1778
rect 3685 -1782 3688 -1778
rect 3674 -1793 3677 -1789
rect 3674 -1813 3677 -1797
rect 3685 -1801 3688 -1789
rect 3685 -1813 3688 -1805
rect 3674 -1825 3677 -1822
rect 3685 -1825 3688 -1822
rect 3678 -1944 3682 -1834
rect 3710 -1851 3714 -1774
rect 3752 -1783 3755 -1779
rect 3763 -1783 3766 -1779
rect 3752 -1794 3755 -1790
rect 3752 -1814 3755 -1798
rect 3763 -1802 3766 -1790
rect 3763 -1814 3766 -1806
rect 3904 -1804 3908 -1705
rect 4015 -1804 4019 -1700
rect 4051 -1725 4055 -1640
rect 4087 -1649 4090 -1645
rect 4098 -1649 4101 -1645
rect 4566 -1655 4569 -1640
rect 4087 -1660 4090 -1656
rect 4087 -1680 4090 -1664
rect 4098 -1668 4101 -1656
rect 4098 -1680 4101 -1672
rect 4566 -1674 4569 -1659
rect 4566 -1683 4569 -1679
rect 4087 -1692 4090 -1689
rect 4098 -1692 4101 -1689
rect 4051 -1728 4073 -1725
rect 4051 -1729 4069 -1728
rect 4066 -1743 4069 -1739
rect 4077 -1743 4080 -1739
rect 4066 -1754 4069 -1750
rect 4066 -1774 4069 -1758
rect 4077 -1762 4080 -1750
rect 4077 -1774 4080 -1766
rect 4066 -1786 4069 -1783
rect 4077 -1786 4080 -1783
rect 4073 -1804 4077 -1795
rect 4094 -1804 4098 -1701
rect 4565 -1804 4569 -1695
rect 5004 -1804 5008 -1069
rect 3904 -1808 5008 -1804
rect 3752 -1826 3755 -1823
rect 3763 -1826 3766 -1823
rect 3710 -1855 3738 -1851
rect 3734 -1862 3738 -1855
rect 3731 -1877 3734 -1873
rect 3742 -1877 3745 -1873
rect 3731 -1888 3734 -1884
rect 3731 -1908 3734 -1892
rect 3742 -1896 3745 -1884
rect 3742 -1908 3745 -1900
rect 3731 -1920 3734 -1917
rect 3742 -1920 3745 -1917
rect 3738 -1944 3742 -1929
rect 3759 -1944 3763 -1835
rect 3904 -1944 3908 -1808
rect 3484 -1948 3908 -1944
<< ndiffusion >>
rect 2985 615 2988 616
rect 2987 611 2988 615
rect 2990 615 2994 616
rect 3004 615 3007 616
rect 2990 611 2992 615
rect 3006 611 3007 615
rect 3009 615 3015 616
rect 3009 611 3011 615
rect 3027 615 3032 616
rect 3031 611 3032 615
rect 3034 615 3037 616
rect 3046 615 3051 616
rect 3034 611 3036 615
rect 3050 611 3051 615
rect 3053 615 3057 616
rect 3053 611 3055 615
rect 3725 631 3728 632
rect 3727 627 3728 631
rect 3730 631 3734 632
rect 3744 631 3747 632
rect 3730 627 3732 631
rect 3746 627 3747 631
rect 3749 631 3755 632
rect 3749 627 3751 631
rect 3767 631 3772 632
rect 3771 627 3772 631
rect 3774 631 3777 632
rect 3786 631 3791 632
rect 3774 627 3776 631
rect 3790 627 3791 631
rect 3793 631 3797 632
rect 3793 627 3795 631
rect 4504 642 4507 643
rect 4506 638 4507 642
rect 4509 642 4513 643
rect 4523 642 4526 643
rect 4509 638 4511 642
rect 4525 638 4526 642
rect 4528 642 4534 643
rect 4528 638 4530 642
rect 4546 642 4551 643
rect 4550 638 4551 642
rect 4553 642 4556 643
rect 4565 642 4570 643
rect 4553 638 4555 642
rect 4569 638 4570 642
rect 4572 642 4576 643
rect 4572 638 4574 642
rect 1263 404 1265 408
rect 1259 399 1265 404
rect 1268 399 1276 408
rect 1279 404 1282 408
rect 1286 404 1287 408
rect 1279 399 1287 404
rect 1086 294 1088 298
rect 1082 289 1088 294
rect 1091 289 1099 298
rect 1102 294 1105 298
rect 1109 294 1110 298
rect 1102 289 1110 294
rect 1143 285 1146 290
rect 1149 285 1153 290
rect 2859 449 2862 450
rect 2861 445 2862 449
rect 2864 449 2868 450
rect 2878 449 2881 450
rect 2864 445 2866 449
rect 2880 445 2881 449
rect 2883 449 2889 450
rect 2883 445 2885 449
rect 2901 449 2906 450
rect 2905 445 2906 449
rect 2908 449 2911 450
rect 2920 449 2925 450
rect 2908 445 2910 449
rect 2924 445 2925 449
rect 2927 449 2931 450
rect 2927 445 2929 449
rect 3064 453 3067 454
rect 3066 449 3067 453
rect 3069 453 3073 454
rect 3083 453 3086 454
rect 3069 449 3071 453
rect 3085 449 3086 453
rect 3088 453 3094 454
rect 3088 449 3090 453
rect 3106 453 3111 454
rect 3110 449 3111 453
rect 3113 453 3116 454
rect 3125 453 3130 454
rect 3113 449 3115 453
rect 3129 449 3130 453
rect 3132 453 3136 454
rect 3132 449 3134 453
rect 1341 403 1343 407
rect 1337 398 1343 403
rect 1346 398 1354 407
rect 1357 403 1360 407
rect 1364 403 1365 407
rect 1357 398 1365 403
rect 1320 309 1322 313
rect 1316 304 1322 309
rect 1325 304 1333 313
rect 1336 309 1339 313
rect 1343 309 1344 313
rect 1336 304 1344 309
rect 1088 211 1090 215
rect 1084 206 1090 211
rect 1093 206 1101 215
rect 1104 211 1107 215
rect 1111 211 1112 215
rect 1104 206 1112 211
rect 1145 202 1148 207
rect 1151 202 1155 207
rect 986 191 989 196
rect 992 191 996 196
rect 987 94 990 99
rect 993 94 997 99
rect 1086 111 1088 115
rect 1082 106 1088 111
rect 1091 106 1099 115
rect 1102 111 1105 115
rect 1109 111 1110 115
rect 1102 106 1110 111
rect 1143 102 1146 107
rect 1149 102 1153 107
rect 1087 22 1089 26
rect 1083 17 1089 22
rect 1092 17 1100 26
rect 1103 22 1106 26
rect 1110 22 1111 26
rect 1103 17 1111 22
rect 1144 13 1147 18
rect 1150 13 1154 18
rect 1427 344 1429 348
rect 1423 339 1429 344
rect 1432 339 1440 348
rect 1443 344 1446 348
rect 1450 344 1451 348
rect 1443 339 1451 344
rect 1538 346 1540 350
rect 1534 341 1540 346
rect 1543 341 1551 350
rect 1554 346 1557 350
rect 1561 346 1562 350
rect 1554 341 1562 346
rect 1654 346 1656 350
rect 1484 335 1487 340
rect 1490 335 1494 340
rect 1595 337 1598 342
rect 1601 337 1605 342
rect 1650 341 1656 346
rect 1659 341 1667 350
rect 1670 346 1673 350
rect 1677 346 1678 350
rect 1670 341 1678 346
rect 1774 347 1776 351
rect 1770 342 1776 347
rect 1779 342 1787 351
rect 1790 347 1793 351
rect 1797 347 1798 351
rect 1790 342 1798 347
rect 1956 348 1958 352
rect 1952 343 1958 348
rect 1961 343 1969 352
rect 1972 348 1975 352
rect 1979 348 1980 352
rect 1972 343 1980 348
rect 2067 350 2069 354
rect 2063 345 2069 350
rect 2072 345 2080 354
rect 2083 350 2086 354
rect 2090 350 2091 354
rect 2083 345 2091 350
rect 2183 350 2185 354
rect 1711 337 1714 342
rect 1717 337 1721 342
rect 1831 338 1834 343
rect 1837 338 1841 343
rect 2013 339 2016 344
rect 2019 339 2023 344
rect 2124 341 2127 346
rect 2130 341 2134 346
rect 2179 345 2185 350
rect 2188 345 2196 354
rect 2199 350 2202 354
rect 2206 350 2207 354
rect 2199 345 2207 350
rect 2303 351 2305 355
rect 2299 346 2305 351
rect 2308 346 2316 355
rect 2319 351 2322 355
rect 2326 351 2327 355
rect 2319 346 2327 351
rect 2860 357 2862 361
rect 2856 352 2862 357
rect 2865 352 2873 361
rect 2876 357 2879 361
rect 2883 357 2884 361
rect 2876 352 2884 357
rect 3015 357 3017 361
rect 2917 348 2920 353
rect 2923 348 2927 353
rect 3011 352 3017 357
rect 3020 352 3028 361
rect 3031 357 3034 361
rect 3038 357 3039 361
rect 3031 352 3039 357
rect 3072 348 3075 353
rect 3078 348 3082 353
rect 2240 341 2243 346
rect 2246 341 2250 346
rect 2360 342 2363 347
rect 2366 342 2370 347
rect 3233 412 3235 416
rect 3229 407 3235 412
rect 3238 407 3246 416
rect 3249 412 3252 416
rect 3256 412 3257 416
rect 3249 407 3257 412
rect 3599 465 3602 466
rect 3601 461 3602 465
rect 3604 465 3608 466
rect 3618 465 3621 466
rect 3604 461 3606 465
rect 3620 461 3621 465
rect 3623 465 3629 466
rect 3623 461 3625 465
rect 3641 465 3646 466
rect 3645 461 3646 465
rect 3648 465 3651 466
rect 3660 465 3665 466
rect 3648 461 3650 465
rect 3664 461 3665 465
rect 3667 465 3671 466
rect 3667 461 3669 465
rect 3804 469 3807 470
rect 3806 465 3807 469
rect 3809 469 3813 470
rect 3823 469 3826 470
rect 3809 465 3811 469
rect 3825 465 3826 469
rect 3828 469 3834 470
rect 3828 465 3830 469
rect 3846 469 3851 470
rect 3850 465 3851 469
rect 3853 469 3856 470
rect 3865 469 3870 470
rect 3853 465 3855 469
rect 3869 465 3870 469
rect 3872 469 3876 470
rect 3872 465 3874 469
rect 5184 636 5187 637
rect 5186 632 5187 636
rect 5189 636 5193 637
rect 5203 636 5206 637
rect 5189 632 5191 636
rect 5205 632 5206 636
rect 5208 636 5214 637
rect 5208 632 5210 636
rect 5226 636 5231 637
rect 5230 632 5231 636
rect 5233 636 5236 637
rect 5245 636 5250 637
rect 5233 632 5235 636
rect 5249 632 5250 636
rect 5252 636 5256 637
rect 5252 632 5254 636
rect 3311 411 3313 415
rect 3307 406 3313 411
rect 3316 406 3324 415
rect 3327 411 3330 415
rect 3334 411 3335 415
rect 3327 406 3335 411
rect 3600 373 3602 377
rect 3596 368 3602 373
rect 3605 368 3613 377
rect 3616 373 3619 377
rect 3623 373 3624 377
rect 3616 368 3624 373
rect 3755 373 3757 377
rect 3657 364 3660 369
rect 3663 364 3667 369
rect 3751 368 3757 373
rect 3760 368 3768 377
rect 3771 373 3774 377
rect 3778 373 3779 377
rect 3771 368 3779 373
rect 3812 364 3815 369
rect 3818 364 3822 369
rect 3973 428 3975 432
rect 3969 423 3975 428
rect 3978 423 3986 432
rect 3989 428 3992 432
rect 3996 428 3997 432
rect 3989 423 3997 428
rect 4378 476 4381 477
rect 4380 472 4381 476
rect 4383 476 4387 477
rect 4397 476 4400 477
rect 4383 472 4385 476
rect 4399 472 4400 476
rect 4402 476 4408 477
rect 4402 472 4404 476
rect 4420 476 4425 477
rect 4424 472 4425 476
rect 4427 476 4430 477
rect 4439 476 4444 477
rect 4427 472 4429 476
rect 4443 472 4444 476
rect 4446 476 4450 477
rect 4446 472 4448 476
rect 4583 480 4586 481
rect 4585 476 4586 480
rect 4588 480 4592 481
rect 4602 480 4605 481
rect 4588 476 4590 480
rect 4604 476 4605 480
rect 4607 480 4613 481
rect 4607 476 4609 480
rect 4625 480 4630 481
rect 4629 476 4630 480
rect 4632 480 4635 481
rect 4644 480 4649 481
rect 4632 476 4634 480
rect 4648 476 4649 480
rect 4651 480 4655 481
rect 4651 476 4653 480
rect 4051 427 4053 431
rect 4047 422 4053 427
rect 4056 422 4064 431
rect 4067 427 4070 431
rect 4074 427 4075 431
rect 4067 422 4075 427
rect 4379 384 4381 388
rect 4375 379 4381 384
rect 4384 379 4392 388
rect 4395 384 4398 388
rect 4402 384 4403 388
rect 4395 379 4403 384
rect 4534 384 4536 388
rect 4436 375 4439 380
rect 4442 375 4446 380
rect 4530 379 4536 384
rect 4539 379 4547 388
rect 4550 384 4553 388
rect 4557 384 4558 388
rect 4550 379 4558 384
rect 4591 375 4594 380
rect 4597 375 4601 380
rect 3290 317 3292 321
rect 3286 312 3292 317
rect 3295 312 3303 321
rect 3306 317 3309 321
rect 3313 317 3314 321
rect 3306 312 3314 317
rect 4030 333 4032 337
rect 4026 328 4032 333
rect 4035 328 4043 337
rect 4046 333 4049 337
rect 4053 333 4054 337
rect 4752 439 4754 443
rect 4748 434 4754 439
rect 4757 434 4765 443
rect 4768 439 4771 443
rect 4775 439 4776 443
rect 4768 434 4776 439
rect 5058 470 5061 471
rect 5060 466 5061 470
rect 5063 470 5067 471
rect 5077 470 5080 471
rect 5063 466 5065 470
rect 5079 466 5080 470
rect 5082 470 5088 471
rect 5082 466 5084 470
rect 5100 470 5105 471
rect 5104 466 5105 470
rect 5107 470 5110 471
rect 5119 470 5124 471
rect 5107 466 5109 470
rect 5123 466 5124 470
rect 5126 470 5130 471
rect 5126 466 5128 470
rect 4830 438 4832 442
rect 4826 433 4832 438
rect 4835 433 4843 442
rect 4846 438 4849 442
rect 4853 438 4854 442
rect 4846 433 4854 438
rect 5263 474 5266 475
rect 5265 470 5266 474
rect 5268 474 5272 475
rect 5282 474 5285 475
rect 5268 470 5270 474
rect 5284 470 5285 474
rect 5287 474 5293 475
rect 5287 470 5289 474
rect 5305 474 5310 475
rect 5309 470 5310 474
rect 5312 474 5315 475
rect 5324 474 5329 475
rect 5312 470 5314 474
rect 5328 470 5329 474
rect 5331 474 5335 475
rect 5331 470 5333 474
rect 5059 378 5061 382
rect 5055 373 5061 378
rect 5064 373 5072 382
rect 5075 378 5078 382
rect 5082 378 5083 382
rect 5075 373 5083 378
rect 5214 378 5216 382
rect 5116 369 5119 374
rect 5122 369 5126 374
rect 5210 373 5216 378
rect 5219 373 5227 382
rect 5230 378 5233 382
rect 5237 378 5238 382
rect 5230 373 5238 378
rect 5271 369 5274 374
rect 5277 369 5281 374
rect 5432 433 5434 437
rect 5428 428 5434 433
rect 5437 428 5445 437
rect 5448 433 5451 437
rect 5455 433 5456 437
rect 5448 428 5456 433
rect 5510 432 5512 436
rect 5506 427 5512 432
rect 5515 427 5523 436
rect 5526 432 5529 436
rect 5533 432 5534 436
rect 5526 427 5534 432
rect 4809 344 4811 348
rect 4805 339 4811 344
rect 4814 339 4822 348
rect 4825 344 4828 348
rect 4832 344 4833 348
rect 4825 339 4833 344
rect 4046 328 4054 333
rect 5489 338 5491 342
rect 5485 333 5491 338
rect 5494 333 5502 342
rect 5505 338 5508 342
rect 5512 338 5513 342
rect 5505 333 5513 338
rect 1430 142 1432 146
rect 1426 137 1432 142
rect 1435 137 1443 146
rect 1446 142 1449 146
rect 1453 142 1454 146
rect 1446 137 1454 142
rect 1541 144 1543 148
rect 1537 139 1543 144
rect 1546 139 1554 148
rect 1557 144 1560 148
rect 1564 144 1565 148
rect 1557 139 1565 144
rect 1657 144 1659 148
rect 1487 133 1490 138
rect 1493 133 1497 138
rect 1598 135 1601 140
rect 1604 135 1608 140
rect 1653 139 1659 144
rect 1662 139 1670 148
rect 1673 144 1676 148
rect 1680 144 1681 148
rect 1673 139 1681 144
rect 1777 145 1779 149
rect 1773 140 1779 145
rect 1782 140 1790 149
rect 1793 145 1796 149
rect 1800 145 1801 149
rect 1793 140 1801 145
rect 1959 146 1961 150
rect 1955 141 1961 146
rect 1964 141 1972 150
rect 1975 146 1978 150
rect 1982 146 1983 150
rect 1975 141 1983 146
rect 2070 148 2072 152
rect 2066 143 2072 148
rect 2075 143 2083 152
rect 2086 148 2089 152
rect 2093 148 2094 152
rect 2086 143 2094 148
rect 2186 148 2188 152
rect 1714 135 1717 140
rect 1720 135 1724 140
rect 1834 136 1837 141
rect 1840 136 1844 141
rect 2016 137 2019 142
rect 2022 137 2026 142
rect 2127 139 2130 144
rect 2133 139 2137 144
rect 2182 143 2188 148
rect 2191 143 2199 152
rect 2202 148 2205 152
rect 2209 148 2210 152
rect 2202 143 2210 148
rect 2306 149 2308 153
rect 2302 144 2308 149
rect 2311 144 2319 153
rect 2322 149 2325 153
rect 2329 149 2330 153
rect 2322 144 2330 149
rect 2243 139 2246 144
rect 2249 139 2253 144
rect 2363 140 2366 145
rect 2369 140 2373 145
rect 1455 -35 1457 -31
rect 1451 -40 1457 -35
rect 1460 -40 1468 -31
rect 1471 -35 1474 -31
rect 1478 -35 1479 -31
rect 1471 -40 1479 -35
rect 1566 -33 1568 -29
rect 1562 -38 1568 -33
rect 1571 -38 1579 -29
rect 1582 -33 1585 -29
rect 1589 -33 1590 -29
rect 1582 -38 1590 -33
rect 1682 -33 1684 -29
rect 1512 -44 1515 -39
rect 1518 -44 1522 -39
rect 1623 -42 1626 -37
rect 1629 -42 1633 -37
rect 1678 -38 1684 -33
rect 1687 -38 1695 -29
rect 1698 -33 1701 -29
rect 1705 -33 1706 -29
rect 1698 -38 1706 -33
rect 1802 -32 1804 -28
rect 1798 -37 1804 -32
rect 1807 -37 1815 -28
rect 1818 -32 1821 -28
rect 1825 -32 1826 -28
rect 1818 -37 1826 -32
rect 1984 -31 1986 -27
rect 1980 -36 1986 -31
rect 1989 -36 1997 -27
rect 2000 -31 2003 -27
rect 2007 -31 2008 -27
rect 2000 -36 2008 -31
rect 2095 -29 2097 -25
rect 2091 -34 2097 -29
rect 2100 -34 2108 -25
rect 2111 -29 2114 -25
rect 2118 -29 2119 -25
rect 2111 -34 2119 -29
rect 2211 -29 2213 -25
rect 1739 -42 1742 -37
rect 1745 -42 1749 -37
rect 1859 -41 1862 -36
rect 1865 -41 1869 -36
rect 2041 -40 2044 -35
rect 2047 -40 2051 -35
rect 2152 -38 2155 -33
rect 2158 -38 2162 -33
rect 2207 -34 2213 -29
rect 2216 -34 2224 -25
rect 2227 -29 2230 -25
rect 2234 -29 2235 -25
rect 2227 -34 2235 -29
rect 2331 -28 2333 -24
rect 2327 -33 2333 -28
rect 2336 -33 2344 -24
rect 2347 -28 2350 -24
rect 2354 -28 2355 -24
rect 2347 -33 2355 -28
rect 2268 -38 2271 -33
rect 2274 -38 2278 -33
rect 2388 -37 2391 -32
rect 2394 -37 2398 -32
rect 1722 -176 1724 -172
rect 1718 -181 1724 -176
rect 1727 -181 1735 -172
rect 1738 -176 1741 -172
rect 1745 -176 1746 -172
rect 1738 -181 1746 -176
rect 1840 -177 1842 -173
rect 1779 -185 1782 -180
rect 1785 -185 1789 -180
rect 1836 -182 1842 -177
rect 1845 -182 1853 -173
rect 1856 -177 1859 -173
rect 1863 -177 1864 -173
rect 1856 -182 1864 -177
rect 1973 -177 1975 -173
rect 1897 -186 1900 -181
rect 1903 -186 1907 -181
rect 1969 -182 1975 -177
rect 1978 -182 1986 -173
rect 1989 -177 1992 -173
rect 1996 -177 1997 -173
rect 1989 -182 1997 -177
rect 2092 -178 2094 -174
rect 2030 -186 2033 -181
rect 2036 -186 2040 -181
rect 2088 -183 2094 -178
rect 2097 -183 2105 -174
rect 2108 -178 2111 -174
rect 2115 -178 2116 -174
rect 2108 -183 2116 -178
rect 2149 -187 2152 -182
rect 2155 -187 2159 -182
rect 3590 -19 3592 -15
rect 3586 -24 3592 -19
rect 3595 -24 3603 -15
rect 3606 -19 3609 -15
rect 3613 -19 3614 -15
rect 3606 -24 3614 -19
rect 3668 -20 3670 -16
rect 3664 -25 3670 -20
rect 3673 -25 3681 -16
rect 3684 -20 3687 -16
rect 3691 -20 3692 -16
rect 3684 -25 3692 -20
rect 3647 -114 3649 -110
rect 3643 -119 3649 -114
rect 3652 -119 3660 -110
rect 3663 -114 3666 -110
rect 3670 -114 3671 -110
rect 3663 -119 3671 -114
rect 3808 -146 3810 -142
rect 3804 -151 3810 -146
rect 3813 -151 3821 -142
rect 3824 -146 3827 -142
rect 3831 -146 3832 -142
rect 3824 -151 3832 -146
rect 3603 -295 3605 -291
rect 3599 -300 3605 -295
rect 3608 -300 3616 -291
rect 3619 -295 3622 -291
rect 3626 -295 3627 -291
rect 3619 -300 3627 -295
rect 3886 -147 3888 -143
rect 3882 -152 3888 -147
rect 3891 -152 3899 -143
rect 3902 -147 3905 -143
rect 3909 -147 3910 -143
rect 3902 -152 3910 -147
rect 3865 -241 3867 -237
rect 3861 -246 3867 -241
rect 3870 -246 3878 -237
rect 3881 -241 3884 -237
rect 3888 -241 3889 -237
rect 3881 -246 3889 -241
rect 4101 -192 4104 -187
rect 4107 -192 4111 -187
rect 3681 -296 3683 -292
rect 3677 -301 3683 -296
rect 3686 -301 3694 -292
rect 3697 -296 3700 -292
rect 3704 -296 3705 -292
rect 3697 -301 3705 -296
rect 3660 -390 3662 -386
rect 3656 -395 3662 -390
rect 3665 -395 3673 -386
rect 3676 -390 3679 -386
rect 3683 -390 3684 -386
rect 3676 -395 3684 -390
rect 2834 -636 2837 -631
rect 2840 -636 2844 -631
rect 2999 -636 3002 -631
rect 3005 -636 3009 -631
rect 3176 -635 3179 -630
rect 3182 -635 3186 -630
rect 3351 -636 3354 -631
rect 3357 -636 3361 -631
rect 3749 -681 3752 -676
rect 3755 -681 3759 -676
rect 2880 -746 2882 -742
rect 2876 -751 2882 -746
rect 2885 -751 2893 -742
rect 2896 -746 2899 -742
rect 2903 -746 2904 -742
rect 2896 -751 2904 -746
rect 3051 -741 3053 -737
rect 3047 -746 3053 -741
rect 3056 -746 3064 -737
rect 3067 -741 3070 -737
rect 3074 -741 3075 -737
rect 3067 -746 3075 -741
rect 3244 -745 3246 -741
rect 3108 -750 3111 -745
rect 3114 -750 3118 -745
rect 3240 -750 3246 -745
rect 3249 -750 3257 -741
rect 3260 -745 3263 -741
rect 3267 -745 3268 -741
rect 3260 -750 3268 -745
rect 3425 -741 3427 -737
rect 3421 -746 3427 -741
rect 3430 -746 3438 -737
rect 3441 -741 3444 -737
rect 3448 -741 3449 -737
rect 3441 -746 3449 -741
rect 2937 -755 2940 -750
rect 2943 -755 2947 -750
rect 3301 -754 3304 -749
rect 3307 -754 3311 -749
rect 3482 -750 3485 -745
rect 3488 -750 3492 -745
rect 3012 -885 3014 -881
rect 3008 -890 3014 -885
rect 3017 -890 3025 -881
rect 3028 -885 3031 -881
rect 3035 -885 3036 -881
rect 3028 -890 3036 -885
rect 3069 -894 3072 -889
rect 3075 -894 3079 -889
rect 3016 -1083 3018 -1079
rect 3012 -1088 3018 -1083
rect 3021 -1088 3029 -1079
rect 3032 -1083 3035 -1079
rect 3039 -1083 3040 -1079
rect 3032 -1088 3040 -1083
rect 3073 -1092 3076 -1087
rect 3079 -1092 3083 -1087
rect 3828 -682 3831 -681
rect 3830 -686 3831 -682
rect 3833 -682 3837 -681
rect 3847 -682 3850 -681
rect 3833 -686 3835 -682
rect 3849 -686 3850 -682
rect 3852 -682 3858 -681
rect 3852 -686 3854 -682
rect 3870 -682 3875 -681
rect 3874 -686 3875 -682
rect 3877 -682 3880 -681
rect 3889 -682 3894 -681
rect 3877 -686 3879 -682
rect 3893 -686 3894 -682
rect 3896 -682 3900 -681
rect 3896 -686 3898 -682
rect 3997 -682 4000 -677
rect 4003 -682 4007 -677
rect 4076 -683 4079 -682
rect 4078 -687 4079 -683
rect 4081 -683 4085 -682
rect 4095 -683 4098 -682
rect 4081 -687 4083 -683
rect 4097 -687 4098 -683
rect 4100 -683 4106 -682
rect 4100 -687 4102 -683
rect 4118 -683 4123 -682
rect 4122 -687 4123 -683
rect 4125 -683 4128 -682
rect 4137 -683 4142 -682
rect 4125 -687 4127 -683
rect 4141 -687 4142 -683
rect 4144 -683 4148 -682
rect 4144 -687 4146 -683
rect 4240 -673 4243 -668
rect 4246 -673 4250 -668
rect 4319 -674 4322 -673
rect 4321 -678 4322 -674
rect 4324 -674 4328 -673
rect 4338 -674 4341 -673
rect 4324 -678 4326 -674
rect 4340 -678 4341 -674
rect 4343 -674 4349 -673
rect 4343 -678 4345 -674
rect 4361 -674 4366 -673
rect 4365 -678 4366 -674
rect 4368 -674 4371 -673
rect 4380 -674 4385 -673
rect 4368 -678 4370 -674
rect 4384 -678 4385 -674
rect 4387 -674 4391 -673
rect 4387 -678 4389 -674
rect 4509 -668 4512 -663
rect 4515 -668 4519 -663
rect 4588 -669 4591 -668
rect 4590 -673 4591 -669
rect 4593 -669 4597 -668
rect 4607 -669 4610 -668
rect 4593 -673 4595 -669
rect 4609 -673 4610 -669
rect 4612 -669 4618 -668
rect 4612 -673 4614 -669
rect 4630 -669 4635 -668
rect 4634 -673 4635 -669
rect 4637 -669 4640 -668
rect 4649 -669 4654 -668
rect 4637 -673 4639 -669
rect 4653 -673 4654 -669
rect 4656 -669 4660 -668
rect 4656 -673 4658 -669
rect 4083 -802 4085 -798
rect 4079 -807 4085 -802
rect 4088 -807 4096 -798
rect 4099 -802 4102 -798
rect 4106 -802 4107 -798
rect 4099 -807 4107 -802
rect 4140 -811 4143 -806
rect 4146 -811 4150 -806
rect 4303 -822 4305 -818
rect 4299 -827 4305 -822
rect 4308 -827 4316 -818
rect 4319 -822 4322 -818
rect 4326 -822 4327 -818
rect 4319 -827 4327 -822
rect 4459 -814 4461 -810
rect 4455 -819 4461 -814
rect 4464 -819 4472 -810
rect 4475 -814 4478 -810
rect 4482 -814 4483 -810
rect 4475 -819 4483 -814
rect 4516 -823 4519 -818
rect 4522 -823 4526 -818
rect 4360 -831 4363 -826
rect 4366 -831 4370 -826
rect 3862 -917 3864 -913
rect 3858 -922 3864 -917
rect 3867 -922 3875 -913
rect 3878 -917 3881 -913
rect 3885 -917 3886 -913
rect 3878 -922 3886 -917
rect 3919 -926 3922 -921
rect 3925 -926 3929 -921
rect 3875 -1103 3877 -1099
rect 3871 -1108 3877 -1103
rect 3880 -1108 3888 -1099
rect 3891 -1103 3894 -1099
rect 3898 -1103 3899 -1099
rect 3891 -1108 3899 -1103
rect 3932 -1112 3935 -1107
rect 3938 -1112 3942 -1107
rect 4203 -1086 4205 -1082
rect 4199 -1091 4205 -1086
rect 4208 -1091 4216 -1082
rect 4219 -1086 4222 -1082
rect 4226 -1086 4227 -1082
rect 4219 -1091 4227 -1086
rect 4260 -1095 4263 -1090
rect 4266 -1095 4270 -1090
rect 2859 -1267 2862 -1262
rect 2865 -1267 2869 -1262
rect 3024 -1267 3027 -1262
rect 3030 -1267 3034 -1262
rect 3201 -1266 3204 -1261
rect 3207 -1266 3211 -1261
rect 3376 -1267 3379 -1262
rect 3382 -1267 3386 -1262
rect 2905 -1377 2907 -1373
rect 2901 -1382 2907 -1377
rect 2910 -1382 2918 -1373
rect 2921 -1377 2924 -1373
rect 2928 -1377 2929 -1373
rect 2921 -1382 2929 -1377
rect 3076 -1372 3078 -1368
rect 3072 -1377 3078 -1372
rect 3081 -1377 3089 -1368
rect 3092 -1372 3095 -1368
rect 3099 -1372 3100 -1368
rect 3092 -1377 3100 -1372
rect 3269 -1376 3271 -1372
rect 3133 -1381 3136 -1376
rect 3139 -1381 3143 -1376
rect 3265 -1381 3271 -1376
rect 3274 -1381 3282 -1372
rect 3285 -1376 3288 -1372
rect 3292 -1376 3293 -1372
rect 3285 -1381 3293 -1376
rect 3450 -1372 3452 -1368
rect 3446 -1377 3452 -1372
rect 3455 -1377 3463 -1368
rect 3466 -1372 3469 -1368
rect 3473 -1372 3474 -1368
rect 3466 -1377 3474 -1372
rect 2962 -1386 2965 -1381
rect 2968 -1386 2972 -1381
rect 3326 -1385 3329 -1380
rect 3332 -1385 3336 -1380
rect 3507 -1381 3510 -1376
rect 3513 -1381 3517 -1376
rect 3662 -1573 3664 -1569
rect 3658 -1578 3664 -1573
rect 3667 -1578 3675 -1569
rect 3678 -1573 3681 -1569
rect 3685 -1573 3686 -1569
rect 3678 -1578 3686 -1573
rect 3740 -1574 3742 -1570
rect 3736 -1579 3742 -1574
rect 3745 -1579 3753 -1570
rect 3756 -1574 3759 -1570
rect 3763 -1574 3764 -1570
rect 3756 -1579 3764 -1574
rect 5013 -1039 5015 -1035
rect 5009 -1044 5015 -1039
rect 5018 -1044 5026 -1035
rect 5029 -1039 5032 -1035
rect 5036 -1039 5037 -1035
rect 5029 -1044 5037 -1039
rect 5230 -1040 5232 -1036
rect 5070 -1048 5073 -1043
rect 5076 -1048 5080 -1043
rect 5226 -1045 5232 -1040
rect 5235 -1045 5243 -1036
rect 5246 -1040 5249 -1036
rect 5253 -1040 5254 -1036
rect 5246 -1045 5254 -1040
rect 5287 -1049 5290 -1044
rect 5293 -1049 5297 -1044
rect 3719 -1668 3721 -1664
rect 3715 -1673 3721 -1668
rect 3724 -1673 3732 -1664
rect 3735 -1668 3738 -1664
rect 3742 -1668 3743 -1664
rect 3735 -1673 3743 -1668
rect 4007 -1683 4009 -1679
rect 4003 -1688 4009 -1683
rect 4012 -1688 4020 -1679
rect 4023 -1683 4026 -1679
rect 4030 -1683 4031 -1679
rect 4023 -1688 4031 -1683
rect 3672 -1817 3674 -1813
rect 3668 -1822 3674 -1817
rect 3677 -1822 3685 -1813
rect 3688 -1817 3691 -1813
rect 3695 -1817 3696 -1813
rect 3688 -1822 3696 -1817
rect 4563 -1679 4566 -1674
rect 4569 -1679 4573 -1674
rect 4085 -1684 4087 -1680
rect 4081 -1689 4087 -1684
rect 4090 -1689 4098 -1680
rect 4101 -1684 4104 -1680
rect 4108 -1684 4109 -1680
rect 4101 -1689 4109 -1684
rect 4064 -1778 4066 -1774
rect 4060 -1783 4066 -1778
rect 4069 -1783 4077 -1774
rect 4080 -1778 4083 -1774
rect 4087 -1778 4088 -1774
rect 4080 -1783 4088 -1778
rect 3750 -1818 3752 -1814
rect 3746 -1823 3752 -1818
rect 3755 -1823 3763 -1814
rect 3766 -1818 3769 -1814
rect 3773 -1818 3774 -1814
rect 3766 -1823 3774 -1818
rect 3729 -1912 3731 -1908
rect 3725 -1917 3731 -1912
rect 3734 -1917 3742 -1908
rect 3745 -1912 3748 -1908
rect 3752 -1912 3753 -1908
rect 3745 -1917 3753 -1912
<< pdiffusion >>
rect 2983 646 2988 647
rect 2987 642 2988 646
rect 2990 646 2996 647
rect 2990 642 2992 646
rect 3002 646 3007 647
rect 3006 642 3007 646
rect 3009 646 3015 647
rect 3009 642 3011 646
rect 3027 646 3032 647
rect 3031 642 3032 646
rect 3034 646 3040 647
rect 3034 642 3036 646
rect 3046 646 3051 647
rect 3050 642 3051 646
rect 3053 646 3059 647
rect 3053 642 3055 646
rect 3723 662 3728 663
rect 3727 658 3728 662
rect 3730 662 3736 663
rect 3730 658 3732 662
rect 3742 662 3747 663
rect 3746 658 3747 662
rect 3749 662 3755 663
rect 3749 658 3751 662
rect 3767 662 3772 663
rect 3771 658 3772 662
rect 3774 662 3780 663
rect 3774 658 3776 662
rect 3786 662 3791 663
rect 3790 658 3791 662
rect 3793 662 3799 663
rect 3793 658 3795 662
rect 4502 673 4507 674
rect 4506 669 4507 673
rect 4509 673 4515 674
rect 4509 669 4511 673
rect 4521 673 4526 674
rect 4525 669 4526 673
rect 4528 673 4534 674
rect 4528 669 4530 673
rect 4546 673 4551 674
rect 4550 669 4551 673
rect 4553 673 4559 674
rect 4553 669 4555 673
rect 4565 673 4570 674
rect 4569 669 4570 673
rect 4572 673 4578 674
rect 4572 669 4574 673
rect 1262 435 1265 439
rect 1258 432 1265 435
rect 1268 435 1271 439
rect 1275 435 1276 439
rect 1268 432 1276 435
rect 1279 435 1282 439
rect 1279 432 1286 435
rect 1085 325 1088 329
rect 1081 322 1088 325
rect 1091 325 1094 329
rect 1098 325 1099 329
rect 1091 322 1099 325
rect 1102 325 1105 329
rect 1102 322 1109 325
rect 1142 324 1146 329
rect 1149 324 1153 329
rect 1157 324 1159 329
rect 1340 434 1343 438
rect 1336 431 1343 434
rect 1346 434 1349 438
rect 1353 434 1354 438
rect 1346 431 1354 434
rect 1357 434 1360 438
rect 1357 431 1364 434
rect 2857 480 2862 481
rect 2861 476 2862 480
rect 2864 480 2870 481
rect 2864 476 2866 480
rect 2876 480 2881 481
rect 2880 476 2881 480
rect 2883 480 2889 481
rect 2883 476 2885 480
rect 2901 480 2906 481
rect 2905 476 2906 480
rect 2908 480 2914 481
rect 2908 476 2910 480
rect 2920 480 2925 481
rect 2924 476 2925 480
rect 2927 480 2933 481
rect 2927 476 2929 480
rect 3062 484 3067 485
rect 3066 480 3067 484
rect 3069 484 3075 485
rect 3069 480 3071 484
rect 3081 484 3086 485
rect 3085 480 3086 484
rect 3088 484 3094 485
rect 3088 480 3090 484
rect 3106 484 3111 485
rect 3110 480 3111 484
rect 3113 484 3119 485
rect 3113 480 3115 484
rect 3125 484 3130 485
rect 3129 480 3130 484
rect 3132 484 3138 485
rect 3132 480 3134 484
rect 3232 443 3235 447
rect 3228 440 3235 443
rect 3238 443 3241 447
rect 3245 443 3246 447
rect 3238 440 3246 443
rect 3249 443 3252 447
rect 3249 440 3256 443
rect 2859 388 2862 392
rect 1319 340 1322 344
rect 1315 337 1322 340
rect 1325 340 1328 344
rect 1332 340 1333 344
rect 1325 337 1333 340
rect 1336 340 1339 344
rect 1336 337 1343 340
rect 1087 242 1090 246
rect 1083 239 1090 242
rect 1093 242 1096 246
rect 1100 242 1101 246
rect 1093 239 1101 242
rect 1104 242 1107 246
rect 1104 239 1111 242
rect 1144 241 1148 246
rect 1151 241 1155 246
rect 1159 241 1161 246
rect 985 230 989 235
rect 992 230 996 235
rect 1000 230 1002 235
rect 986 133 990 138
rect 993 133 997 138
rect 1001 133 1003 138
rect 1085 142 1088 146
rect 1081 139 1088 142
rect 1091 142 1094 146
rect 1098 142 1099 146
rect 1091 139 1099 142
rect 1102 142 1105 146
rect 1102 139 1109 142
rect 1142 141 1146 146
rect 1149 141 1153 146
rect 1157 141 1159 146
rect 1086 53 1089 57
rect 1082 50 1089 53
rect 1092 53 1095 57
rect 1099 53 1100 57
rect 1092 50 1100 53
rect 1103 53 1106 57
rect 1103 50 1110 53
rect 1143 52 1147 57
rect 1150 52 1154 57
rect 1158 52 1160 57
rect 1426 375 1429 379
rect 1422 372 1429 375
rect 1432 375 1435 379
rect 1439 375 1440 379
rect 1432 372 1440 375
rect 1443 375 1446 379
rect 1443 372 1450 375
rect 1483 374 1487 379
rect 1490 374 1494 379
rect 1498 374 1500 379
rect 1537 377 1540 381
rect 1533 374 1540 377
rect 1543 377 1546 381
rect 1550 377 1551 381
rect 1543 374 1551 377
rect 1554 377 1557 381
rect 1554 374 1561 377
rect 1594 376 1598 381
rect 1601 376 1605 381
rect 1609 376 1611 381
rect 1653 377 1656 381
rect 1649 374 1656 377
rect 1659 377 1662 381
rect 1666 377 1667 381
rect 1659 374 1667 377
rect 1670 377 1673 381
rect 1670 374 1677 377
rect 1710 376 1714 381
rect 1717 376 1721 381
rect 1725 376 1727 381
rect 1773 378 1776 382
rect 1769 375 1776 378
rect 1779 378 1782 382
rect 1786 378 1787 382
rect 1779 375 1787 378
rect 1790 378 1793 382
rect 1790 375 1797 378
rect 1830 377 1834 382
rect 1837 377 1841 382
rect 1845 377 1847 382
rect 1955 379 1958 383
rect 1951 376 1958 379
rect 1961 379 1964 383
rect 1968 379 1969 383
rect 1961 376 1969 379
rect 1972 379 1975 383
rect 1972 376 1979 379
rect 2012 378 2016 383
rect 2019 378 2023 383
rect 2027 378 2029 383
rect 2066 381 2069 385
rect 2062 378 2069 381
rect 2072 381 2075 385
rect 2079 381 2080 385
rect 2072 378 2080 381
rect 2083 381 2086 385
rect 2083 378 2090 381
rect 2123 380 2127 385
rect 2130 380 2134 385
rect 2138 380 2140 385
rect 2182 381 2185 385
rect 2178 378 2185 381
rect 2188 381 2191 385
rect 2195 381 2196 385
rect 2188 378 2196 381
rect 2199 381 2202 385
rect 2199 378 2206 381
rect 2239 380 2243 385
rect 2246 380 2250 385
rect 2254 380 2256 385
rect 2302 382 2305 386
rect 2298 379 2305 382
rect 2308 382 2311 386
rect 2315 382 2316 386
rect 2308 379 2316 382
rect 2319 382 2322 386
rect 2319 379 2326 382
rect 2359 381 2363 386
rect 2366 381 2370 386
rect 2374 381 2376 386
rect 2855 385 2862 388
rect 2865 388 2868 392
rect 2872 388 2873 392
rect 2865 385 2873 388
rect 2876 388 2879 392
rect 2876 385 2883 388
rect 2916 387 2920 392
rect 2923 387 2927 392
rect 2931 387 2933 392
rect 3014 388 3017 392
rect 3010 385 3017 388
rect 3020 388 3023 392
rect 3027 388 3028 392
rect 3020 385 3028 388
rect 3031 388 3034 392
rect 3031 385 3038 388
rect 3071 387 3075 392
rect 3078 387 3082 392
rect 3086 387 3088 392
rect 3597 496 3602 497
rect 3601 492 3602 496
rect 3604 496 3610 497
rect 3604 492 3606 496
rect 3616 496 3621 497
rect 3620 492 3621 496
rect 3623 496 3629 497
rect 3623 492 3625 496
rect 3641 496 3646 497
rect 3645 492 3646 496
rect 3648 496 3654 497
rect 3648 492 3650 496
rect 3660 496 3665 497
rect 3664 492 3665 496
rect 3667 496 3673 497
rect 3667 492 3669 496
rect 3310 442 3313 446
rect 3306 439 3313 442
rect 3316 442 3319 446
rect 3323 442 3324 446
rect 3316 439 3324 442
rect 3327 442 3330 446
rect 3327 439 3334 442
rect 3802 500 3807 501
rect 3806 496 3807 500
rect 3809 500 3815 501
rect 3809 496 3811 500
rect 3821 500 3826 501
rect 3825 496 3826 500
rect 3828 500 3834 501
rect 3828 496 3830 500
rect 3846 500 3851 501
rect 3850 496 3851 500
rect 3853 500 3859 501
rect 3853 496 3855 500
rect 3865 500 3870 501
rect 3869 496 3870 500
rect 3872 500 3878 501
rect 3872 496 3874 500
rect 5182 667 5187 668
rect 5186 663 5187 667
rect 5189 667 5195 668
rect 5189 663 5191 667
rect 5201 667 5206 668
rect 5205 663 5206 667
rect 5208 667 5214 668
rect 5208 663 5210 667
rect 5226 667 5231 668
rect 5230 663 5231 667
rect 5233 667 5239 668
rect 5233 663 5235 667
rect 5245 667 5250 668
rect 5249 663 5250 667
rect 5252 667 5258 668
rect 5252 663 5254 667
rect 3972 459 3975 463
rect 3968 456 3975 459
rect 3978 459 3981 463
rect 3985 459 3986 463
rect 3978 456 3986 459
rect 3989 459 3992 463
rect 3989 456 3996 459
rect 3599 404 3602 408
rect 3595 401 3602 404
rect 3605 404 3608 408
rect 3612 404 3613 408
rect 3605 401 3613 404
rect 3616 404 3619 408
rect 3616 401 3623 404
rect 3656 403 3660 408
rect 3663 403 3667 408
rect 3671 403 3673 408
rect 3754 404 3757 408
rect 3750 401 3757 404
rect 3760 404 3763 408
rect 3767 404 3768 408
rect 3760 401 3768 404
rect 3771 404 3774 408
rect 3771 401 3778 404
rect 3811 403 3815 408
rect 3818 403 3822 408
rect 3826 403 3828 408
rect 3289 348 3292 352
rect 3285 345 3292 348
rect 3295 348 3298 352
rect 3302 348 3303 352
rect 3295 345 3303 348
rect 3306 348 3309 352
rect 3306 345 3313 348
rect 4050 458 4053 462
rect 4046 455 4053 458
rect 4056 458 4059 462
rect 4063 458 4064 462
rect 4056 455 4064 458
rect 4067 458 4070 462
rect 4376 507 4381 508
rect 4380 503 4381 507
rect 4383 507 4389 508
rect 4383 503 4385 507
rect 4395 507 4400 508
rect 4399 503 4400 507
rect 4402 507 4408 508
rect 4402 503 4404 507
rect 4420 507 4425 508
rect 4424 503 4425 507
rect 4427 507 4433 508
rect 4427 503 4429 507
rect 4439 507 4444 508
rect 4443 503 4444 507
rect 4446 507 4452 508
rect 4446 503 4448 507
rect 4067 455 4074 458
rect 4581 511 4586 512
rect 4585 507 4586 511
rect 4588 511 4594 512
rect 4588 507 4590 511
rect 4600 511 4605 512
rect 4604 507 4605 511
rect 4607 511 4613 512
rect 4607 507 4609 511
rect 4625 511 4630 512
rect 4629 507 4630 511
rect 4632 511 4638 512
rect 4632 507 4634 511
rect 4644 511 4649 512
rect 4648 507 4649 511
rect 4651 511 4657 512
rect 4651 507 4653 511
rect 4751 470 4754 474
rect 4747 467 4754 470
rect 4757 470 4760 474
rect 4764 470 4765 474
rect 4757 467 4765 470
rect 4768 470 4771 474
rect 4768 467 4775 470
rect 4378 415 4381 419
rect 4374 412 4381 415
rect 4384 415 4387 419
rect 4391 415 4392 419
rect 4384 412 4392 415
rect 4395 415 4398 419
rect 4395 412 4402 415
rect 4435 414 4439 419
rect 4442 414 4446 419
rect 4450 414 4452 419
rect 4533 415 4536 419
rect 4529 412 4536 415
rect 4539 415 4542 419
rect 4546 415 4547 419
rect 4539 412 4547 415
rect 4550 415 4553 419
rect 4550 412 4557 415
rect 4590 414 4594 419
rect 4597 414 4601 419
rect 4605 414 4607 419
rect 4029 364 4032 368
rect 4025 361 4032 364
rect 4035 364 4038 368
rect 4042 364 4043 368
rect 4035 361 4043 364
rect 4046 364 4049 368
rect 4046 361 4053 364
rect 4829 469 4832 473
rect 4825 466 4832 469
rect 4835 469 4838 473
rect 4842 469 4843 473
rect 4835 466 4843 469
rect 4846 469 4849 473
rect 4846 466 4853 469
rect 5056 501 5061 502
rect 5060 497 5061 501
rect 5063 501 5069 502
rect 5063 497 5065 501
rect 5075 501 5080 502
rect 5079 497 5080 501
rect 5082 501 5088 502
rect 5082 497 5084 501
rect 5100 501 5105 502
rect 5104 497 5105 501
rect 5107 501 5113 502
rect 5107 497 5109 501
rect 5119 501 5124 502
rect 5123 497 5124 501
rect 5126 501 5132 502
rect 5126 497 5128 501
rect 5261 505 5266 506
rect 5265 501 5266 505
rect 5268 505 5274 506
rect 5268 501 5270 505
rect 5280 505 5285 506
rect 5284 501 5285 505
rect 5287 505 5293 506
rect 5287 501 5289 505
rect 5305 505 5310 506
rect 5309 501 5310 505
rect 5312 505 5318 506
rect 5312 501 5314 505
rect 5324 505 5329 506
rect 5328 501 5329 505
rect 5331 505 5337 506
rect 5331 501 5333 505
rect 5431 464 5434 468
rect 5427 461 5434 464
rect 5437 464 5440 468
rect 5444 464 5445 468
rect 5437 461 5445 464
rect 5448 464 5451 468
rect 5448 461 5455 464
rect 5058 409 5061 413
rect 5054 406 5061 409
rect 5064 409 5067 413
rect 5071 409 5072 413
rect 5064 406 5072 409
rect 5075 409 5078 413
rect 5075 406 5082 409
rect 5115 408 5119 413
rect 5122 408 5126 413
rect 5130 408 5132 413
rect 5213 409 5216 413
rect 5209 406 5216 409
rect 5219 409 5222 413
rect 5226 409 5227 413
rect 5219 406 5227 409
rect 5230 409 5233 413
rect 5230 406 5237 409
rect 5270 408 5274 413
rect 5277 408 5281 413
rect 5285 408 5287 413
rect 4808 375 4811 379
rect 4804 372 4811 375
rect 4814 375 4817 379
rect 4821 375 4822 379
rect 4814 372 4822 375
rect 4825 375 4828 379
rect 4825 372 4832 375
rect 5509 463 5512 467
rect 5505 460 5512 463
rect 5515 463 5518 467
rect 5522 463 5523 467
rect 5515 460 5523 463
rect 5526 463 5529 467
rect 5526 460 5533 463
rect 5488 369 5491 373
rect 5484 366 5491 369
rect 5494 369 5497 373
rect 5501 369 5502 373
rect 5494 366 5502 369
rect 5505 369 5508 373
rect 5505 366 5512 369
rect 1429 173 1432 177
rect 1425 170 1432 173
rect 1435 173 1438 177
rect 1442 173 1443 177
rect 1435 170 1443 173
rect 1446 173 1449 177
rect 1446 170 1453 173
rect 1486 172 1490 177
rect 1493 172 1497 177
rect 1501 172 1503 177
rect 1540 175 1543 179
rect 1536 172 1543 175
rect 1546 175 1549 179
rect 1553 175 1554 179
rect 1546 172 1554 175
rect 1557 175 1560 179
rect 1557 172 1564 175
rect 1597 174 1601 179
rect 1604 174 1608 179
rect 1612 174 1614 179
rect 1656 175 1659 179
rect 1652 172 1659 175
rect 1662 175 1665 179
rect 1669 175 1670 179
rect 1662 172 1670 175
rect 1673 175 1676 179
rect 1673 172 1680 175
rect 1713 174 1717 179
rect 1720 174 1724 179
rect 1728 174 1730 179
rect 1776 176 1779 180
rect 1772 173 1779 176
rect 1782 176 1785 180
rect 1789 176 1790 180
rect 1782 173 1790 176
rect 1793 176 1796 180
rect 1793 173 1800 176
rect 1833 175 1837 180
rect 1840 175 1844 180
rect 1848 175 1850 180
rect 1958 177 1961 181
rect 1954 174 1961 177
rect 1964 177 1967 181
rect 1971 177 1972 181
rect 1964 174 1972 177
rect 1975 177 1978 181
rect 1975 174 1982 177
rect 2015 176 2019 181
rect 2022 176 2026 181
rect 2030 176 2032 181
rect 2069 179 2072 183
rect 2065 176 2072 179
rect 2075 179 2078 183
rect 2082 179 2083 183
rect 2075 176 2083 179
rect 2086 179 2089 183
rect 2086 176 2093 179
rect 2126 178 2130 183
rect 2133 178 2137 183
rect 2141 178 2143 183
rect 2185 179 2188 183
rect 2181 176 2188 179
rect 2191 179 2194 183
rect 2198 179 2199 183
rect 2191 176 2199 179
rect 2202 179 2205 183
rect 2202 176 2209 179
rect 2242 178 2246 183
rect 2249 178 2253 183
rect 2257 178 2259 183
rect 2305 180 2308 184
rect 2301 177 2308 180
rect 2311 180 2314 184
rect 2318 180 2319 184
rect 2311 177 2319 180
rect 2322 180 2325 184
rect 2322 177 2329 180
rect 2362 179 2366 184
rect 2369 179 2373 184
rect 2377 179 2379 184
rect 1454 -2 1457 1
rect 1450 -5 1457 -2
rect 1460 -2 1463 1
rect 1467 -2 1468 1
rect 1460 -5 1468 -2
rect 1471 -2 1474 1
rect 1471 -5 1478 -2
rect 1511 -3 1515 1
rect 1518 -3 1522 1
rect 1526 -3 1528 1
rect 1565 -2 1568 1
rect 1561 -5 1568 -2
rect 1571 -2 1574 1
rect 1578 -2 1579 1
rect 1571 -5 1579 -2
rect 1582 -2 1585 1
rect 1582 -5 1589 -2
rect 1622 -3 1626 1
rect 1629 -3 1633 1
rect 1637 -3 1639 1
rect 1681 -2 1684 1
rect 1687 -2 1690 1
rect 1694 -2 1695 1
rect 1698 -2 1701 1
rect 1738 -4 1742 0
rect 1745 -4 1749 0
rect 1753 -4 1755 0
rect 1801 -1 1804 2
rect 1807 -1 1810 2
rect 1814 -1 1815 2
rect 1818 -1 1821 2
rect 1983 1 1986 4
rect 1989 1 1992 4
rect 1996 1 1997 4
rect 2000 1 2003 4
rect 1858 -4 1862 0
rect 1865 -4 1869 0
rect 1873 -4 1875 0
rect 2040 0 2044 4
rect 2047 0 2051 4
rect 2055 0 2057 4
rect 2094 3 2097 6
rect 2100 3 2103 6
rect 2107 3 2108 6
rect 2111 3 2114 6
rect 2151 3 2155 6
rect 2158 3 2162 6
rect 2166 3 2168 6
rect 2210 3 2213 6
rect 2216 3 2219 6
rect 2223 3 2224 6
rect 2227 3 2230 6
rect 2267 3 2271 6
rect 2274 3 2278 6
rect 2282 3 2284 6
rect 2330 3 2333 7
rect 2336 3 2339 7
rect 2343 3 2344 7
rect 2347 3 2350 7
rect 2387 3 2391 7
rect 2394 3 2398 7
rect 2402 3 2404 7
rect 1721 -145 1724 -141
rect 1717 -148 1724 -145
rect 1727 -145 1730 -141
rect 1734 -145 1735 -141
rect 1727 -148 1735 -145
rect 1738 -145 1741 -141
rect 1738 -148 1745 -145
rect 1778 -146 1782 -141
rect 1785 -146 1789 -141
rect 1793 -146 1795 -141
rect 1839 -146 1842 -142
rect 1835 -149 1842 -146
rect 1845 -146 1848 -142
rect 1852 -146 1853 -142
rect 1845 -149 1853 -146
rect 1856 -146 1859 -142
rect 1856 -149 1863 -146
rect 1896 -147 1900 -142
rect 1903 -147 1907 -142
rect 1911 -147 1913 -142
rect 1972 -146 1975 -142
rect 1968 -149 1975 -146
rect 1978 -146 1981 -142
rect 1985 -146 1986 -142
rect 1978 -149 1986 -146
rect 1989 -146 1992 -142
rect 1989 -149 1996 -146
rect 2029 -147 2033 -142
rect 2036 -147 2040 -142
rect 2044 -147 2046 -142
rect 2091 -147 2094 -143
rect 2087 -150 2094 -147
rect 2097 -147 2100 -143
rect 2104 -147 2105 -143
rect 2097 -150 2105 -147
rect 2108 -147 2111 -143
rect 2108 -150 2115 -147
rect 2148 -148 2152 -143
rect 2155 -148 2159 -143
rect 2163 -148 2165 -143
rect 3589 12 3592 16
rect 3585 9 3592 12
rect 3595 12 3598 16
rect 3602 12 3603 16
rect 3595 9 3603 12
rect 3606 12 3609 16
rect 3606 9 3613 12
rect 3667 11 3670 15
rect 3663 8 3670 11
rect 3673 11 3676 15
rect 3680 11 3681 15
rect 3673 8 3681 11
rect 3684 11 3687 15
rect 3684 8 3691 11
rect 3646 -83 3649 -79
rect 3642 -86 3649 -83
rect 3652 -83 3655 -79
rect 3659 -83 3660 -79
rect 3652 -86 3660 -83
rect 3663 -83 3666 -79
rect 3663 -86 3670 -83
rect 3807 -115 3810 -111
rect 3803 -118 3810 -115
rect 3813 -115 3816 -111
rect 3820 -115 3821 -111
rect 3813 -118 3821 -115
rect 3824 -115 3827 -111
rect 3824 -118 3831 -115
rect 3885 -116 3888 -112
rect 3881 -119 3888 -116
rect 3891 -116 3894 -112
rect 3898 -116 3899 -112
rect 3891 -119 3899 -116
rect 3902 -116 3905 -112
rect 3902 -119 3909 -116
rect 3602 -264 3605 -260
rect 3598 -267 3605 -264
rect 3608 -264 3611 -260
rect 3615 -264 3616 -260
rect 3608 -267 3616 -264
rect 3619 -264 3622 -260
rect 3619 -267 3626 -264
rect 3680 -265 3683 -261
rect 3676 -268 3683 -265
rect 3686 -265 3689 -261
rect 3693 -265 3694 -261
rect 3686 -268 3694 -265
rect 3697 -265 3700 -261
rect 3697 -268 3704 -265
rect 4100 -153 4104 -148
rect 4107 -153 4111 -148
rect 4115 -153 4117 -148
rect 3864 -210 3867 -206
rect 3860 -213 3867 -210
rect 3870 -210 3873 -206
rect 3877 -210 3878 -206
rect 3870 -213 3878 -210
rect 3881 -210 3884 -206
rect 3881 -213 3888 -210
rect 3659 -359 3662 -355
rect 3655 -362 3662 -359
rect 3665 -359 3668 -355
rect 3672 -359 3673 -355
rect 3665 -362 3673 -359
rect 3676 -359 3679 -355
rect 3676 -362 3683 -359
rect 2833 -597 2837 -592
rect 2840 -597 2844 -592
rect 2848 -597 2850 -592
rect 2998 -597 3002 -592
rect 3005 -597 3009 -592
rect 3013 -597 3015 -592
rect 3175 -596 3179 -591
rect 3182 -596 3186 -591
rect 3190 -596 3192 -591
rect 3350 -597 3354 -592
rect 3357 -597 3361 -592
rect 3365 -597 3367 -592
rect 3748 -642 3752 -637
rect 3755 -642 3759 -637
rect 3763 -642 3765 -637
rect 3050 -710 3053 -706
rect 2879 -715 2882 -711
rect 2875 -718 2882 -715
rect 2885 -715 2888 -711
rect 2892 -715 2893 -711
rect 2885 -718 2893 -715
rect 2896 -715 2899 -711
rect 2896 -718 2903 -715
rect 2936 -716 2940 -711
rect 2943 -716 2947 -711
rect 2951 -716 2953 -711
rect 3046 -713 3053 -710
rect 3056 -710 3059 -706
rect 3063 -710 3064 -706
rect 3056 -713 3064 -710
rect 3067 -710 3070 -706
rect 3067 -713 3074 -710
rect 3107 -711 3111 -706
rect 3114 -711 3118 -706
rect 3122 -711 3124 -706
rect 3424 -710 3427 -706
rect 3243 -714 3246 -710
rect 3239 -717 3246 -714
rect 3249 -714 3252 -710
rect 3256 -714 3257 -710
rect 3249 -717 3257 -714
rect 3260 -714 3263 -710
rect 3260 -717 3267 -714
rect 3300 -715 3304 -710
rect 3307 -715 3311 -710
rect 3315 -715 3317 -710
rect 3420 -713 3427 -710
rect 3430 -710 3433 -706
rect 3437 -710 3438 -706
rect 3430 -713 3438 -710
rect 3441 -710 3444 -706
rect 3441 -713 3448 -710
rect 3481 -711 3485 -706
rect 3488 -711 3492 -706
rect 3496 -711 3498 -706
rect 3011 -854 3014 -850
rect 3007 -857 3014 -854
rect 3017 -854 3020 -850
rect 3024 -854 3025 -850
rect 3017 -857 3025 -854
rect 3028 -854 3031 -850
rect 3028 -857 3035 -854
rect 3068 -855 3072 -850
rect 3075 -855 3079 -850
rect 3083 -855 3085 -850
rect 3015 -1052 3018 -1048
rect 3011 -1055 3018 -1052
rect 3021 -1052 3024 -1048
rect 3028 -1052 3029 -1048
rect 3021 -1055 3029 -1052
rect 3032 -1052 3035 -1048
rect 3032 -1055 3039 -1052
rect 3072 -1053 3076 -1048
rect 3079 -1053 3083 -1048
rect 3087 -1053 3089 -1048
rect 3996 -643 4000 -638
rect 4003 -643 4007 -638
rect 4011 -643 4013 -638
rect 3826 -651 3831 -650
rect 3830 -655 3831 -651
rect 3833 -651 3839 -650
rect 3833 -655 3835 -651
rect 3845 -651 3850 -650
rect 3849 -655 3850 -651
rect 3852 -651 3858 -650
rect 3852 -655 3854 -651
rect 3870 -651 3875 -650
rect 3874 -655 3875 -651
rect 3877 -651 3883 -650
rect 3877 -655 3879 -651
rect 3889 -651 3894 -650
rect 3893 -655 3894 -651
rect 3896 -651 3902 -650
rect 3896 -655 3898 -651
rect 4239 -634 4243 -629
rect 4246 -634 4250 -629
rect 4254 -634 4256 -629
rect 4074 -652 4079 -651
rect 4078 -656 4079 -652
rect 4081 -652 4087 -651
rect 4081 -656 4083 -652
rect 4093 -652 4098 -651
rect 4097 -656 4098 -652
rect 4100 -652 4106 -651
rect 4100 -656 4102 -652
rect 4118 -652 4123 -651
rect 4122 -656 4123 -652
rect 4125 -652 4131 -651
rect 4125 -656 4127 -652
rect 4137 -652 4142 -651
rect 4141 -656 4142 -652
rect 4144 -652 4150 -651
rect 4144 -656 4146 -652
rect 4508 -629 4512 -624
rect 4515 -629 4519 -624
rect 4523 -629 4525 -624
rect 4317 -643 4322 -642
rect 4321 -647 4322 -643
rect 4324 -643 4330 -642
rect 4324 -647 4326 -643
rect 4336 -643 4341 -642
rect 4340 -647 4341 -643
rect 4343 -643 4349 -642
rect 4343 -647 4345 -643
rect 4361 -643 4366 -642
rect 4365 -647 4366 -643
rect 4368 -643 4374 -642
rect 4368 -647 4370 -643
rect 4380 -643 4385 -642
rect 4384 -647 4385 -643
rect 4387 -643 4393 -642
rect 4387 -647 4389 -643
rect 4586 -638 4591 -637
rect 4590 -642 4591 -638
rect 4593 -638 4599 -637
rect 4593 -642 4595 -638
rect 4605 -638 4610 -637
rect 4609 -642 4610 -638
rect 4612 -638 4618 -637
rect 4612 -642 4614 -638
rect 4630 -638 4635 -637
rect 4634 -642 4635 -638
rect 4637 -638 4643 -637
rect 4637 -642 4639 -638
rect 4649 -638 4654 -637
rect 4653 -642 4654 -638
rect 4656 -638 4662 -637
rect 4656 -642 4658 -638
rect 4082 -771 4085 -767
rect 4078 -774 4085 -771
rect 4088 -771 4091 -767
rect 4095 -771 4096 -767
rect 4088 -774 4096 -771
rect 4099 -771 4102 -767
rect 4099 -774 4106 -771
rect 4139 -772 4143 -767
rect 4146 -772 4150 -767
rect 4154 -772 4156 -767
rect 4458 -783 4461 -779
rect 4454 -786 4461 -783
rect 4464 -783 4467 -779
rect 4471 -783 4472 -779
rect 4464 -786 4472 -783
rect 4475 -783 4478 -779
rect 4475 -786 4482 -783
rect 4515 -784 4519 -779
rect 4522 -784 4526 -779
rect 4530 -784 4532 -779
rect 4302 -791 4305 -787
rect 4298 -794 4305 -791
rect 4308 -791 4311 -787
rect 4315 -791 4316 -787
rect 4308 -794 4316 -791
rect 4319 -791 4322 -787
rect 4319 -794 4326 -791
rect 4359 -792 4363 -787
rect 4366 -792 4370 -787
rect 4374 -792 4376 -787
rect 3861 -886 3864 -882
rect 3857 -889 3864 -886
rect 3867 -886 3870 -882
rect 3874 -886 3875 -882
rect 3867 -889 3875 -886
rect 3878 -886 3881 -882
rect 3878 -889 3885 -886
rect 3918 -887 3922 -882
rect 3925 -887 3929 -882
rect 3933 -887 3935 -882
rect 3874 -1072 3877 -1068
rect 3870 -1075 3877 -1072
rect 3880 -1072 3883 -1068
rect 3887 -1072 3888 -1068
rect 3880 -1075 3888 -1072
rect 3891 -1072 3894 -1068
rect 3891 -1075 3898 -1072
rect 3931 -1073 3935 -1068
rect 3938 -1073 3942 -1068
rect 3946 -1073 3948 -1068
rect 4202 -1055 4205 -1051
rect 4198 -1058 4205 -1055
rect 4208 -1055 4211 -1051
rect 4215 -1055 4216 -1051
rect 4208 -1058 4216 -1055
rect 4219 -1055 4222 -1051
rect 4219 -1058 4226 -1055
rect 4259 -1056 4263 -1051
rect 4266 -1056 4270 -1051
rect 4274 -1056 4276 -1051
rect 2858 -1228 2862 -1223
rect 2865 -1228 2869 -1223
rect 2873 -1228 2875 -1223
rect 3023 -1228 3027 -1223
rect 3030 -1228 3034 -1223
rect 3038 -1228 3040 -1223
rect 3200 -1227 3204 -1222
rect 3207 -1227 3211 -1222
rect 3215 -1227 3217 -1222
rect 3375 -1228 3379 -1223
rect 3382 -1228 3386 -1223
rect 3390 -1228 3392 -1223
rect 3075 -1341 3078 -1337
rect 2904 -1346 2907 -1342
rect 2900 -1349 2907 -1346
rect 2910 -1346 2913 -1342
rect 2917 -1346 2918 -1342
rect 2910 -1349 2918 -1346
rect 2921 -1346 2924 -1342
rect 2921 -1349 2928 -1346
rect 2961 -1347 2965 -1342
rect 2968 -1347 2972 -1342
rect 2976 -1347 2978 -1342
rect 3071 -1344 3078 -1341
rect 3081 -1341 3084 -1337
rect 3088 -1341 3089 -1337
rect 3081 -1344 3089 -1341
rect 3092 -1341 3095 -1337
rect 3092 -1344 3099 -1341
rect 3132 -1342 3136 -1337
rect 3139 -1342 3143 -1337
rect 3147 -1342 3149 -1337
rect 3449 -1341 3452 -1337
rect 3268 -1345 3271 -1341
rect 3264 -1348 3271 -1345
rect 3274 -1345 3277 -1341
rect 3281 -1345 3282 -1341
rect 3274 -1348 3282 -1345
rect 3285 -1345 3288 -1341
rect 3285 -1348 3292 -1345
rect 3325 -1346 3329 -1341
rect 3332 -1346 3336 -1341
rect 3340 -1346 3342 -1341
rect 3445 -1344 3452 -1341
rect 3455 -1341 3458 -1337
rect 3462 -1341 3463 -1337
rect 3455 -1344 3463 -1341
rect 3466 -1341 3469 -1337
rect 3466 -1344 3473 -1341
rect 3506 -1342 3510 -1337
rect 3513 -1342 3517 -1337
rect 3521 -1342 3523 -1337
rect 3661 -1542 3664 -1538
rect 3657 -1545 3664 -1542
rect 3667 -1542 3670 -1538
rect 3674 -1542 3675 -1538
rect 3667 -1545 3675 -1542
rect 3678 -1542 3681 -1538
rect 3678 -1545 3685 -1542
rect 3739 -1543 3742 -1539
rect 3735 -1546 3742 -1543
rect 3745 -1543 3748 -1539
rect 3752 -1543 3753 -1539
rect 3745 -1546 3753 -1543
rect 3756 -1543 3759 -1539
rect 3756 -1546 3763 -1543
rect 5012 -1008 5015 -1004
rect 5008 -1011 5015 -1008
rect 5018 -1008 5021 -1004
rect 5025 -1008 5026 -1004
rect 5018 -1011 5026 -1008
rect 5029 -1008 5032 -1004
rect 5029 -1011 5036 -1008
rect 5069 -1009 5073 -1004
rect 5076 -1009 5080 -1004
rect 5084 -1009 5086 -1004
rect 5229 -1009 5232 -1005
rect 5225 -1012 5232 -1009
rect 5235 -1009 5238 -1005
rect 5242 -1009 5243 -1005
rect 5235 -1012 5243 -1009
rect 5246 -1009 5249 -1005
rect 5246 -1012 5253 -1009
rect 5286 -1010 5290 -1005
rect 5293 -1010 5297 -1005
rect 5301 -1010 5303 -1005
rect 3718 -1637 3721 -1633
rect 3714 -1640 3721 -1637
rect 3724 -1637 3727 -1633
rect 3731 -1637 3732 -1633
rect 3724 -1640 3732 -1637
rect 3735 -1637 3738 -1633
rect 3735 -1640 3742 -1637
rect 4562 -1640 4566 -1635
rect 4569 -1640 4573 -1635
rect 4577 -1640 4579 -1635
rect 4006 -1652 4009 -1648
rect 4002 -1655 4009 -1652
rect 4012 -1652 4015 -1648
rect 4019 -1652 4020 -1648
rect 4012 -1655 4020 -1652
rect 4023 -1652 4026 -1648
rect 4023 -1655 4030 -1652
rect 3671 -1786 3674 -1782
rect 3667 -1789 3674 -1786
rect 3677 -1786 3680 -1782
rect 3684 -1786 3685 -1782
rect 3677 -1789 3685 -1786
rect 3688 -1786 3691 -1782
rect 3688 -1789 3695 -1786
rect 3749 -1787 3752 -1783
rect 3745 -1790 3752 -1787
rect 3755 -1787 3758 -1783
rect 3762 -1787 3763 -1783
rect 3755 -1790 3763 -1787
rect 3766 -1787 3769 -1783
rect 3766 -1790 3773 -1787
rect 4084 -1653 4087 -1649
rect 4080 -1656 4087 -1653
rect 4090 -1653 4093 -1649
rect 4097 -1653 4098 -1649
rect 4090 -1656 4098 -1653
rect 4101 -1653 4104 -1649
rect 4101 -1656 4108 -1653
rect 4063 -1747 4066 -1743
rect 4059 -1750 4066 -1747
rect 4069 -1747 4072 -1743
rect 4076 -1747 4077 -1743
rect 4069 -1750 4077 -1747
rect 4080 -1747 4083 -1743
rect 4080 -1750 4087 -1747
rect 3728 -1881 3731 -1877
rect 3724 -1884 3731 -1881
rect 3734 -1881 3737 -1877
rect 3741 -1881 3742 -1877
rect 3734 -1884 3742 -1881
rect 3745 -1881 3748 -1877
rect 3745 -1884 3752 -1881
<< metal1 >>
rect 741 990 5799 1013
rect 741 988 3035 990
rect 741 263 766 988
rect 3039 988 3776 990
rect 3780 988 4555 990
rect 4559 988 5233 990
rect 5237 988 5799 990
rect 4104 771 4257 775
rect 3364 755 3439 759
rect 2755 701 3015 704
rect 1258 447 1297 448
rect 1301 447 1364 448
rect 1258 445 1316 447
rect 1258 439 1262 445
rect 1282 439 1286 445
rect 1320 445 1364 447
rect 1336 444 1364 445
rect 1336 438 1340 444
rect 1360 438 1364 444
rect 1271 428 1275 435
rect 1215 424 1264 428
rect 1271 425 1286 428
rect 1349 427 1353 434
rect 1081 337 1118 339
rect 1122 337 1141 339
rect 1081 335 1141 337
rect 1145 335 1170 339
rect 1081 329 1085 335
rect 1105 329 1109 335
rect 1138 329 1141 335
rect 1094 318 1098 325
rect 1042 314 1087 318
rect 1094 315 1109 318
rect 741 259 764 263
rect 741 154 766 259
rect 971 241 984 245
rect 988 243 991 245
rect 995 243 1012 245
rect 988 241 1012 243
rect 981 235 984 241
rect 968 211 988 215
rect 997 213 1000 230
rect 1042 213 1046 314
rect 1105 312 1109 315
rect 997 208 1046 213
rect 997 196 1000 208
rect 981 184 985 191
rect 971 180 1013 184
rect 971 178 987 180
rect 991 178 1013 180
rect 741 150 764 154
rect 741 37 766 150
rect 972 144 985 148
rect 989 144 993 148
rect 997 144 1013 148
rect 982 138 985 144
rect 998 118 1001 133
rect 1042 135 1046 208
rect 1062 306 1098 310
rect 1105 309 1110 312
rect 1154 310 1157 324
rect 1215 310 1219 424
rect 1257 420 1260 424
rect 1282 422 1286 425
rect 1332 423 1342 427
rect 1349 424 1364 427
rect 1257 416 1275 420
rect 1282 419 1287 422
rect 1334 419 1338 423
rect 1360 421 1364 424
rect 1360 419 1365 421
rect 1282 415 1294 419
rect 1334 415 1353 419
rect 1360 416 1372 419
rect 1282 408 1286 415
rect 1259 395 1263 404
rect 1259 393 1288 395
rect 1259 392 1271 393
rect 1275 392 1281 393
rect 1285 392 1288 393
rect 1291 325 1294 415
rect 1360 407 1364 416
rect 1337 394 1341 403
rect 1337 391 1366 394
rect 1352 389 1354 391
rect 1369 365 1372 416
rect 1936 403 2283 407
rect 1407 402 2283 403
rect 1407 398 1941 402
rect 1407 382 1412 398
rect 1297 362 1372 365
rect 1384 378 1412 382
rect 1297 333 1301 362
rect 1315 352 1316 354
rect 1325 354 1332 357
rect 1320 352 1343 354
rect 1315 350 1343 352
rect 1315 344 1319 350
rect 1339 344 1343 350
rect 1328 333 1332 340
rect 1297 329 1321 333
rect 1328 330 1343 333
rect 1339 327 1343 330
rect 1384 327 1388 378
rect 1407 368 1412 378
rect 1422 385 1458 389
rect 1462 385 1482 389
rect 1486 385 1511 389
rect 1422 379 1426 385
rect 1446 379 1450 385
rect 1479 379 1482 385
rect 1435 368 1439 375
rect 1407 364 1428 368
rect 1435 365 1450 368
rect 1421 356 1439 360
rect 1446 359 1450 365
rect 1495 359 1498 374
rect 1517 370 1522 398
rect 1533 388 1570 391
rect 1574 388 1593 391
rect 1533 387 1593 388
rect 1597 387 1622 391
rect 1533 381 1537 387
rect 1557 381 1561 387
rect 1590 381 1593 387
rect 1546 370 1550 377
rect 1517 366 1539 370
rect 1546 367 1561 370
rect 1557 364 1561 367
rect 1446 355 1486 359
rect 1495 356 1505 359
rect 1532 358 1550 362
rect 1557 361 1562 364
rect 1606 361 1609 376
rect 1635 370 1640 398
rect 1649 389 1685 391
rect 1689 389 1709 391
rect 1649 387 1709 389
rect 1713 387 1738 391
rect 1649 381 1653 387
rect 1673 381 1677 387
rect 1706 381 1709 387
rect 1662 370 1666 377
rect 1635 366 1655 370
rect 1662 367 1677 370
rect 1673 364 1677 367
rect 1446 348 1450 355
rect 1423 335 1427 344
rect 1495 340 1498 356
rect 1423 332 1469 335
rect 1479 332 1483 335
rect 1451 331 1483 332
rect 1451 329 1461 331
rect 1465 329 1483 331
rect 1291 321 1332 325
rect 1339 323 1388 327
rect 1339 313 1343 323
rect 1062 227 1066 306
rect 1105 305 1145 309
rect 1154 306 1219 310
rect 1105 298 1109 305
rect 1082 285 1086 294
rect 1154 290 1157 306
rect 1316 300 1320 309
rect 1316 297 1345 300
rect 1327 296 1335 297
rect 1327 295 1328 296
rect 1332 295 1335 296
rect 1082 283 1128 285
rect 1138 283 1142 285
rect 1082 282 1142 283
rect 1110 280 1142 282
rect 1138 279 1142 280
rect 1138 275 1140 279
rect 1368 275 1391 280
rect 1083 254 1121 256
rect 1125 254 1143 256
rect 1083 252 1143 254
rect 1147 252 1172 256
rect 1083 246 1087 252
rect 1107 246 1111 252
rect 1140 246 1143 252
rect 1096 235 1100 242
rect 1081 231 1089 235
rect 1096 232 1111 235
rect 1107 229 1111 232
rect 1062 223 1100 227
rect 1107 226 1112 229
rect 1156 226 1159 241
rect 1042 131 1044 135
rect 1062 118 1066 223
rect 1107 222 1147 226
rect 1156 222 1160 226
rect 1107 215 1111 222
rect 1084 202 1088 211
rect 1156 207 1159 222
rect 1502 216 1505 356
rect 1557 357 1597 361
rect 1606 358 1621 361
rect 1648 358 1666 362
rect 1673 361 1678 364
rect 1557 350 1561 357
rect 1534 337 1538 346
rect 1606 342 1609 358
rect 1534 334 1580 337
rect 1590 334 1594 337
rect 1562 333 1594 334
rect 1562 331 1572 333
rect 1576 331 1594 333
rect 1618 247 1621 358
rect 1673 357 1713 361
rect 1722 360 1725 376
rect 1749 371 1754 398
rect 1769 390 1807 392
rect 1811 390 1829 392
rect 1769 388 1829 390
rect 1833 388 1858 392
rect 1769 382 1773 388
rect 1793 382 1797 388
rect 1826 382 1829 388
rect 1782 371 1786 378
rect 1749 367 1775 371
rect 1782 368 1797 371
rect 1793 365 1797 368
rect 1722 357 1741 360
rect 1769 359 1786 363
rect 1793 362 1798 365
rect 1673 350 1677 357
rect 1650 337 1654 346
rect 1722 342 1725 357
rect 1650 334 1696 337
rect 1706 334 1710 337
rect 1678 333 1710 334
rect 1678 331 1686 333
rect 1690 331 1710 333
rect 1738 257 1741 357
rect 1793 358 1833 362
rect 1842 360 1845 377
rect 1935 372 1941 398
rect 1951 391 1989 393
rect 1993 391 2011 393
rect 1951 389 2011 391
rect 2015 389 2040 393
rect 1951 383 1955 389
rect 1975 383 1979 389
rect 2008 383 2011 389
rect 1964 372 1968 379
rect 1935 368 1957 372
rect 1964 369 1979 372
rect 1950 360 1968 364
rect 1975 363 1979 369
rect 2024 363 2027 378
rect 2046 374 2051 402
rect 2062 393 2101 395
rect 2105 393 2122 395
rect 2062 391 2122 393
rect 2126 391 2151 395
rect 2062 385 2066 391
rect 2086 385 2090 391
rect 2119 385 2122 391
rect 2075 374 2079 381
rect 2046 370 2068 374
rect 2075 371 2090 374
rect 2086 368 2090 371
rect 1793 351 1797 358
rect 1842 356 1896 360
rect 1770 338 1774 347
rect 1842 343 1845 356
rect 1770 335 1816 338
rect 1826 335 1830 338
rect 1798 334 1830 335
rect 1798 332 1808 334
rect 1812 332 1830 334
rect 1892 323 1896 356
rect 1975 359 2015 363
rect 2024 359 2026 363
rect 2061 362 2079 366
rect 2086 365 2091 368
rect 2135 366 2138 380
rect 2164 374 2169 402
rect 2178 393 2217 395
rect 2221 393 2238 395
rect 2178 391 2238 393
rect 2242 391 2267 395
rect 2178 385 2182 391
rect 2202 385 2206 391
rect 2235 385 2238 391
rect 2191 374 2195 381
rect 2164 370 2184 374
rect 2191 371 2206 374
rect 2202 368 2206 371
rect 2086 361 2126 365
rect 2135 362 2137 366
rect 2177 362 2195 366
rect 2202 365 2207 368
rect 1975 352 1979 359
rect 1952 339 1956 348
rect 2024 344 2027 359
rect 2086 354 2090 361
rect 2063 341 2067 350
rect 2135 346 2138 362
rect 2202 361 2242 365
rect 2251 364 2254 380
rect 2278 375 2283 402
rect 2298 394 2335 396
rect 2339 394 2358 396
rect 2298 392 2358 394
rect 2362 392 2387 396
rect 2298 386 2302 392
rect 2322 386 2326 392
rect 2355 386 2358 392
rect 2311 375 2315 382
rect 2278 371 2304 375
rect 2311 372 2326 375
rect 2322 369 2326 372
rect 2202 354 2206 361
rect 2251 360 2252 364
rect 2294 363 2296 367
rect 2300 363 2315 367
rect 2322 366 2327 369
rect 2322 362 2362 366
rect 2371 362 2374 381
rect 2755 362 2758 701
rect 3010 674 3015 701
rect 2983 670 3023 674
rect 2983 646 2987 670
rect 2983 615 2987 642
rect 2992 646 2996 667
rect 3000 663 3015 667
rect 3011 646 3015 663
rect 2992 615 2996 642
rect 3002 615 3006 642
rect 3011 615 3015 642
rect 3019 630 3023 670
rect 3027 660 3035 662
rect 3039 660 3050 662
rect 3027 658 3050 660
rect 3027 646 3031 658
rect 3046 646 3050 658
rect 3019 626 3029 630
rect 3036 622 3040 642
rect 3055 630 3059 642
rect 3047 626 3048 630
rect 3055 626 3058 630
rect 3019 618 3040 622
rect 3002 608 3006 611
rect 3019 608 3023 618
rect 3036 615 3040 618
rect 3055 615 3059 626
rect 3002 604 3023 608
rect 3027 608 3031 611
rect 3046 609 3050 611
rect 3045 608 3050 609
rect 3027 604 3050 608
rect 2179 341 2183 350
rect 2251 346 2254 360
rect 2322 355 2326 362
rect 2371 359 2758 362
rect 2782 523 2892 527
rect 2782 381 2786 523
rect 2888 508 2892 523
rect 2857 504 2897 508
rect 2857 480 2861 504
rect 2857 449 2861 476
rect 2866 497 2885 501
rect 2866 480 2870 497
rect 2885 480 2889 497
rect 2866 449 2870 476
rect 2876 449 2880 476
rect 2885 449 2889 476
rect 2893 465 2897 504
rect 2901 494 2916 496
rect 2920 494 2924 496
rect 2901 492 2924 494
rect 2901 480 2905 492
rect 2920 480 2924 492
rect 2893 464 2898 465
rect 2893 460 2903 464
rect 2910 456 2914 476
rect 2929 464 2933 476
rect 2919 457 2922 463
rect 2929 460 2932 464
rect 2893 452 2914 456
rect 2876 442 2880 445
rect 2893 442 2897 452
rect 2910 449 2914 452
rect 2929 449 2933 460
rect 2876 438 2897 442
rect 2901 442 2905 445
rect 2918 443 2924 445
rect 2917 442 2924 443
rect 2901 438 2924 442
rect 2920 425 2924 438
rect 3031 425 3035 604
rect 3062 508 3092 512
rect 3096 508 3102 512
rect 3062 484 3066 508
rect 3062 453 3066 480
rect 3071 501 3094 505
rect 3071 484 3075 501
rect 3090 484 3094 501
rect 3071 453 3075 480
rect 3081 453 3085 480
rect 3090 453 3094 480
rect 3098 468 3102 508
rect 3106 498 3113 500
rect 3117 501 3119 502
rect 3117 500 3122 501
rect 3117 498 3129 500
rect 3106 496 3129 498
rect 3106 484 3110 496
rect 3125 484 3129 496
rect 3098 464 3108 468
rect 3115 460 3119 480
rect 3134 468 3138 480
rect 3123 461 3127 468
rect 3134 464 3137 468
rect 3098 456 3119 460
rect 3126 457 3127 461
rect 3081 446 3085 449
rect 3098 446 3102 456
rect 3115 453 3119 456
rect 3134 453 3138 464
rect 3238 457 3250 458
rect 3081 442 3102 446
rect 3228 455 3274 457
rect 3278 456 3321 457
rect 3278 455 3334 456
rect 3228 453 3334 455
rect 3106 446 3110 449
rect 3125 448 3129 449
rect 3122 446 3129 448
rect 3106 445 3129 446
rect 3105 442 3129 445
rect 3228 447 3232 453
rect 3252 447 3256 453
rect 3306 452 3334 453
rect 3306 446 3310 452
rect 3330 446 3334 452
rect 3107 425 3111 442
rect 3241 436 3245 443
rect 2920 423 3111 425
rect 2920 421 3103 423
rect 3107 421 3111 423
rect 3202 432 3234 436
rect 3241 433 3256 436
rect 3319 435 3323 442
rect 2855 400 2892 402
rect 3020 402 3032 403
rect 2896 400 2915 402
rect 2855 398 2915 400
rect 2919 398 2944 402
rect 3010 400 3047 402
rect 3051 400 3070 402
rect 3010 398 3070 400
rect 3074 398 3099 402
rect 2855 392 2859 398
rect 2879 392 2883 398
rect 2912 392 2915 398
rect 3010 392 3014 398
rect 3034 392 3038 398
rect 2868 381 2872 388
rect 3067 392 3070 398
rect 2782 377 2861 381
rect 2868 378 2883 381
rect 2299 342 2303 351
rect 2371 347 2374 359
rect 1952 336 1998 339
rect 2008 336 2012 339
rect 2063 338 2109 341
rect 2119 338 2123 341
rect 2179 338 2225 341
rect 2235 338 2239 341
rect 2299 339 2345 342
rect 2355 339 2359 342
rect 1980 335 2012 336
rect 2091 337 2123 338
rect 2091 335 2101 337
rect 1980 333 1990 335
rect 1994 333 2012 335
rect 2105 335 2123 337
rect 2207 337 2239 338
rect 2207 335 2217 337
rect 2221 335 2239 337
rect 2327 338 2359 339
rect 2327 336 2337 338
rect 2341 336 2359 338
rect 2782 323 2786 377
rect 2879 375 2883 378
rect 2854 369 2872 373
rect 2879 372 2884 375
rect 2928 372 2931 387
rect 3023 381 3027 388
rect 3009 377 3016 381
rect 3023 378 3038 381
rect 3034 375 3038 378
rect 2879 368 2919 372
rect 2928 369 2954 372
rect 3008 369 3027 373
rect 3034 372 3039 375
rect 3083 373 3086 387
rect 2879 361 2883 368
rect 2856 348 2860 357
rect 2928 353 2931 369
rect 2856 347 2888 348
rect 2912 347 2916 348
rect 2856 346 2916 347
rect 2856 345 2888 346
rect 2884 344 2888 345
rect 2892 344 2916 346
rect 1892 319 2786 323
rect 2951 321 2954 369
rect 3034 368 3074 372
rect 3083 369 3088 373
rect 3034 361 3038 368
rect 3011 348 3015 357
rect 3083 353 3086 369
rect 3011 345 3057 348
rect 3038 344 3058 345
rect 3067 344 3071 348
rect 3038 343 3071 344
rect 3039 341 3046 343
rect 3051 341 3071 343
rect 3202 321 3205 432
rect 3227 428 3230 432
rect 3252 430 3256 433
rect 3304 431 3312 435
rect 3319 432 3334 435
rect 3227 424 3245 428
rect 3252 427 3257 430
rect 3304 427 3308 431
rect 3330 429 3334 432
rect 3330 427 3335 429
rect 3252 423 3264 427
rect 3304 423 3323 427
rect 3330 424 3342 427
rect 3252 416 3256 423
rect 3229 403 3233 412
rect 3229 400 3258 403
rect 3229 345 3233 400
rect 3236 398 3239 400
rect 3243 398 3246 400
rect 3231 341 3233 345
rect 2951 318 3205 321
rect 3229 301 3233 341
rect 3261 333 3264 423
rect 3330 415 3334 424
rect 3307 402 3311 411
rect 3307 400 3336 402
rect 3307 399 3318 400
rect 3316 397 3318 399
rect 3322 399 3336 400
rect 3322 397 3324 399
rect 3339 373 3342 424
rect 3267 370 3342 373
rect 3267 341 3271 370
rect 3292 363 3294 365
rect 3298 363 3303 365
rect 3292 362 3303 363
rect 3285 358 3313 362
rect 3285 352 3289 358
rect 3309 352 3313 358
rect 3298 341 3302 348
rect 3267 337 3291 341
rect 3298 338 3313 341
rect 3309 335 3313 338
rect 3261 329 3302 333
rect 3309 332 3326 335
rect 3309 331 3321 332
rect 3309 321 3313 331
rect 3286 308 3290 317
rect 3286 305 3315 308
rect 3300 301 3304 305
rect 3229 297 3304 301
rect 3434 262 3438 755
rect 3723 688 3753 690
rect 3757 688 3763 690
rect 3723 686 3763 688
rect 3723 662 3727 686
rect 3723 631 3727 658
rect 3732 662 3736 683
rect 3740 679 3755 683
rect 3751 662 3755 679
rect 3732 631 3736 658
rect 3742 631 3746 658
rect 3751 631 3755 658
rect 3759 646 3763 686
rect 3767 676 3776 678
rect 3780 676 3790 678
rect 3767 674 3790 676
rect 3767 662 3771 674
rect 3786 662 3790 674
rect 3759 642 3769 646
rect 3776 638 3780 658
rect 3795 646 3799 658
rect 3787 642 3788 646
rect 3795 642 3798 646
rect 3759 634 3780 638
rect 3742 624 3746 627
rect 3759 624 3763 634
rect 3776 631 3780 634
rect 3795 631 3799 642
rect 3742 620 3763 624
rect 3767 624 3771 627
rect 3786 625 3790 627
rect 3785 624 3790 625
rect 3767 620 3790 624
rect 3574 534 3632 538
rect 3574 397 3578 534
rect 3628 524 3632 534
rect 3597 520 3637 524
rect 3597 496 3601 520
rect 3597 465 3601 492
rect 3606 513 3625 517
rect 3606 512 3611 513
rect 3606 496 3610 512
rect 3625 496 3629 513
rect 3606 465 3610 492
rect 3616 465 3620 492
rect 3625 465 3629 492
rect 3633 481 3637 520
rect 3641 509 3651 512
rect 3655 509 3664 512
rect 3641 508 3664 509
rect 3641 496 3645 508
rect 3660 496 3664 508
rect 3633 480 3638 481
rect 3633 476 3643 480
rect 3650 472 3654 492
rect 3669 480 3673 492
rect 3659 473 3662 479
rect 3669 476 3672 480
rect 3633 468 3654 472
rect 3616 458 3620 461
rect 3633 458 3637 468
rect 3650 465 3654 468
rect 3669 465 3673 476
rect 3616 454 3637 458
rect 3641 458 3645 461
rect 3658 459 3664 461
rect 3657 458 3664 459
rect 3641 454 3664 458
rect 3648 446 3652 454
rect 3767 446 3771 620
rect 3802 524 3832 528
rect 3836 524 3842 528
rect 3802 500 3806 524
rect 3802 469 3806 496
rect 3811 517 3834 521
rect 3811 500 3815 517
rect 3830 500 3834 517
rect 3811 469 3815 496
rect 3821 469 3825 496
rect 3830 469 3834 496
rect 3838 484 3842 524
rect 3846 514 3856 516
rect 3860 514 3869 516
rect 3846 512 3869 514
rect 3846 500 3850 512
rect 3865 500 3869 512
rect 3838 480 3848 484
rect 3855 476 3859 496
rect 3874 484 3878 496
rect 3863 477 3867 484
rect 3874 480 3877 484
rect 3838 472 3859 476
rect 3866 473 3867 477
rect 3821 462 3825 465
rect 3838 462 3842 472
rect 3855 469 3859 472
rect 3874 469 3878 480
rect 3978 473 3990 474
rect 3821 458 3842 462
rect 3968 471 4020 473
rect 4024 472 4061 473
rect 4024 471 4074 472
rect 3968 469 4074 471
rect 3846 462 3850 465
rect 3865 464 3869 465
rect 3862 462 3869 464
rect 3846 461 3869 462
rect 3845 458 3869 461
rect 3968 463 3972 469
rect 3992 463 3996 469
rect 4046 468 4074 469
rect 4046 462 4050 468
rect 4070 462 4074 468
rect 3853 446 3857 458
rect 3981 452 3985 459
rect 3648 444 3857 446
rect 3648 442 3849 444
rect 3853 442 3857 444
rect 3942 448 3974 452
rect 3981 449 3996 452
rect 4059 451 4063 458
rect 3595 416 3629 418
rect 3760 418 3772 419
rect 3633 416 3655 418
rect 3595 414 3655 416
rect 3659 414 3684 418
rect 3750 416 3787 418
rect 3791 416 3810 418
rect 3750 414 3810 416
rect 3814 414 3839 418
rect 3595 408 3599 414
rect 3619 408 3623 414
rect 3652 408 3655 414
rect 3750 408 3754 414
rect 3774 408 3778 414
rect 3608 397 3612 404
rect 3807 408 3810 414
rect 3556 393 3601 397
rect 3608 394 3623 397
rect 3619 391 3623 394
rect 3594 385 3612 389
rect 3619 388 3624 391
rect 3668 388 3671 403
rect 3763 397 3767 404
rect 3749 393 3756 397
rect 3763 394 3778 397
rect 3774 391 3778 394
rect 3619 384 3659 388
rect 3668 385 3694 388
rect 3748 385 3767 389
rect 3774 388 3779 391
rect 3823 389 3826 403
rect 3619 377 3623 384
rect 3596 364 3600 373
rect 3668 369 3671 385
rect 3596 363 3628 364
rect 3652 363 3656 364
rect 3596 362 3656 363
rect 3596 361 3635 362
rect 3624 360 3635 361
rect 3639 360 3656 362
rect 3691 337 3694 385
rect 3774 384 3814 388
rect 3823 385 3828 389
rect 3774 377 3778 384
rect 3751 364 3755 373
rect 3823 369 3826 385
rect 3751 361 3797 364
rect 3778 360 3798 361
rect 3807 360 3811 364
rect 3778 359 3811 360
rect 3779 358 3811 359
rect 3779 356 3791 358
rect 3795 357 3811 358
rect 3795 356 3839 357
rect 3803 351 3839 356
rect 3942 337 3945 448
rect 3967 444 3970 448
rect 3992 446 3996 449
rect 4044 447 4052 451
rect 4059 448 4074 451
rect 3967 440 3985 444
rect 3992 443 3997 446
rect 4044 443 4048 447
rect 4070 445 4074 448
rect 4070 443 4075 445
rect 3992 439 4004 443
rect 4044 439 4063 443
rect 4070 440 4082 443
rect 3992 432 3996 439
rect 3969 419 3973 428
rect 3969 417 3998 419
rect 3969 416 3970 417
rect 3974 416 3998 417
rect 3974 414 3986 416
rect 4001 349 4004 439
rect 4070 431 4074 440
rect 4047 418 4051 427
rect 4047 416 4076 418
rect 4049 415 4076 416
rect 4049 412 4064 415
rect 4079 389 4082 440
rect 4007 386 4082 389
rect 4007 357 4011 386
rect 4032 379 4038 381
rect 4042 379 4043 381
rect 4032 378 4043 379
rect 4025 374 4053 378
rect 4025 368 4029 374
rect 4049 368 4053 374
rect 4038 357 4042 364
rect 4007 353 4031 357
rect 4038 354 4053 357
rect 4049 351 4053 354
rect 4001 345 4042 349
rect 4049 347 4074 351
rect 4049 337 4053 347
rect 3691 334 3945 337
rect 4026 325 4030 333
rect 4028 324 4030 325
rect 4028 321 4055 324
rect 4037 319 4048 321
rect 4070 262 4074 347
rect 4253 289 4257 771
rect 5240 743 5243 833
rect 5161 740 5243 743
rect 4502 698 4534 701
rect 4538 698 4542 701
rect 4502 697 4542 698
rect 4502 673 4506 697
rect 4502 642 4506 669
rect 4511 673 4515 694
rect 4519 690 4534 694
rect 4530 673 4534 690
rect 4511 642 4515 669
rect 4521 642 4525 669
rect 4530 642 4534 669
rect 4538 657 4542 697
rect 4546 687 4555 689
rect 4559 687 4569 689
rect 4546 685 4569 687
rect 4546 673 4550 685
rect 4565 673 4569 685
rect 4538 653 4548 657
rect 4555 649 4559 669
rect 4574 657 4578 669
rect 4566 653 4567 657
rect 4574 653 4577 657
rect 4538 645 4559 649
rect 4521 635 4525 638
rect 4538 635 4542 645
rect 4555 642 4559 645
rect 4574 642 4578 653
rect 4521 631 4542 635
rect 4546 635 4550 638
rect 4565 636 4569 638
rect 4564 635 4569 636
rect 4546 631 4569 635
rect 4357 543 4411 546
rect 4357 408 4361 543
rect 4407 535 4411 543
rect 4376 531 4416 535
rect 4376 507 4380 531
rect 4376 476 4380 503
rect 4385 524 4404 528
rect 4385 523 4390 524
rect 4385 507 4389 523
rect 4404 507 4408 524
rect 4385 476 4389 503
rect 4395 476 4399 503
rect 4404 476 4408 503
rect 4412 492 4416 531
rect 4420 521 4428 523
rect 4432 521 4443 523
rect 4420 519 4443 521
rect 4420 507 4424 519
rect 4439 507 4443 519
rect 4412 491 4417 492
rect 4412 487 4422 491
rect 4429 483 4433 503
rect 4448 491 4452 503
rect 4438 484 4441 490
rect 4448 487 4451 491
rect 4412 479 4433 483
rect 4395 469 4399 472
rect 4412 469 4416 479
rect 4429 476 4433 479
rect 4448 476 4452 487
rect 4395 465 4416 469
rect 4420 469 4424 472
rect 4437 470 4443 472
rect 4436 469 4443 470
rect 4420 465 4443 469
rect 4420 455 4424 465
rect 4547 455 4551 631
rect 5037 543 5091 546
rect 4581 535 4611 539
rect 4615 535 4621 539
rect 4581 511 4585 535
rect 4581 480 4585 507
rect 4590 528 4613 532
rect 4590 511 4594 528
rect 4609 511 4613 528
rect 4590 480 4594 507
rect 4600 480 4604 507
rect 4609 480 4613 507
rect 4617 495 4621 535
rect 4625 525 4633 527
rect 4637 525 4648 527
rect 4625 523 4648 525
rect 4625 511 4629 523
rect 4644 511 4648 523
rect 4617 491 4627 495
rect 4634 487 4638 507
rect 4653 495 4657 507
rect 4642 488 4646 495
rect 4653 491 4656 495
rect 4617 483 4638 487
rect 4645 484 4646 488
rect 4600 473 4604 476
rect 4617 473 4621 483
rect 4634 480 4638 483
rect 4653 480 4657 491
rect 4757 484 4769 485
rect 4600 469 4621 473
rect 4747 482 4789 484
rect 4794 483 4840 484
rect 4794 482 4853 483
rect 4747 480 4853 482
rect 4625 473 4629 476
rect 4644 475 4648 476
rect 4641 473 4648 475
rect 4625 472 4648 473
rect 4624 469 4648 472
rect 4747 474 4751 480
rect 4771 474 4775 480
rect 4825 479 4853 480
rect 4825 473 4829 479
rect 4849 473 4853 479
rect 4629 455 4633 469
rect 4760 463 4764 470
rect 4420 453 4633 455
rect 4420 451 4627 453
rect 4631 451 4633 453
rect 4721 459 4753 463
rect 4760 460 4775 463
rect 4838 462 4842 469
rect 4374 427 4409 429
rect 4539 429 4551 430
rect 4413 427 4434 429
rect 4374 425 4434 427
rect 4438 425 4463 429
rect 4529 427 4566 429
rect 4570 427 4589 429
rect 4529 425 4589 427
rect 4593 425 4618 429
rect 4374 419 4378 425
rect 4398 419 4402 425
rect 4431 419 4434 425
rect 4529 419 4533 425
rect 4553 419 4557 425
rect 4387 408 4391 415
rect 4586 419 4589 425
rect 4335 404 4380 408
rect 4387 405 4402 408
rect 4398 402 4402 405
rect 4373 396 4391 400
rect 4398 399 4403 402
rect 4447 399 4450 414
rect 4542 408 4546 415
rect 4528 404 4535 408
rect 4542 405 4557 408
rect 4553 402 4557 405
rect 4398 395 4438 399
rect 4447 396 4473 399
rect 4527 396 4546 400
rect 4553 399 4558 402
rect 4602 400 4605 414
rect 4398 388 4402 395
rect 4375 375 4379 384
rect 4447 380 4450 396
rect 4375 374 4407 375
rect 4431 374 4435 375
rect 4375 373 4435 374
rect 4375 372 4411 373
rect 4403 371 4411 372
rect 4415 371 4435 373
rect 4470 348 4473 396
rect 4553 395 4593 399
rect 4602 396 4607 400
rect 4553 388 4557 395
rect 4530 375 4534 384
rect 4602 380 4605 396
rect 4530 372 4576 375
rect 4557 371 4577 372
rect 4586 371 4590 375
rect 4557 370 4590 371
rect 4558 369 4590 370
rect 4558 367 4565 369
rect 4569 368 4590 369
rect 4569 367 4618 368
rect 4576 362 4618 367
rect 4721 348 4724 459
rect 4746 455 4749 459
rect 4771 457 4775 460
rect 4823 458 4831 462
rect 4838 459 4853 462
rect 4746 451 4764 455
rect 4771 454 4776 457
rect 4823 454 4827 458
rect 4849 456 4853 459
rect 4849 454 4854 456
rect 4771 450 4783 454
rect 4823 450 4842 454
rect 4849 451 4861 454
rect 4771 443 4775 450
rect 4748 430 4752 439
rect 4748 428 4777 430
rect 4748 427 4750 428
rect 4754 427 4777 428
rect 4757 425 4758 427
rect 4762 425 4765 427
rect 4780 360 4783 450
rect 4849 442 4853 451
rect 4826 429 4830 438
rect 4826 426 4855 429
rect 4835 424 4837 426
rect 4841 424 4843 426
rect 4858 400 4861 451
rect 4786 397 4861 400
rect 5037 402 5040 543
rect 5087 529 5091 543
rect 5056 525 5096 529
rect 5056 501 5060 525
rect 5056 470 5060 497
rect 5065 518 5084 522
rect 5065 517 5070 518
rect 5065 501 5069 517
rect 5084 501 5088 518
rect 5065 470 5069 497
rect 5075 470 5079 497
rect 5084 470 5088 497
rect 5092 486 5096 525
rect 5100 515 5110 517
rect 5114 515 5123 517
rect 5100 513 5123 515
rect 5100 501 5104 513
rect 5119 501 5123 513
rect 5092 485 5097 486
rect 5092 481 5102 485
rect 5109 477 5113 497
rect 5128 485 5132 497
rect 5118 478 5121 484
rect 5128 481 5131 485
rect 5092 473 5113 477
rect 5075 463 5079 466
rect 5092 463 5096 473
rect 5109 470 5113 473
rect 5128 470 5132 481
rect 5075 459 5096 463
rect 5100 463 5104 466
rect 5117 464 5123 466
rect 5116 463 5123 464
rect 5100 459 5123 463
rect 5108 450 5112 459
rect 5108 445 5152 450
rect 5054 421 5089 423
rect 5094 421 5114 423
rect 5054 419 5114 421
rect 5118 419 5143 423
rect 5054 413 5058 419
rect 5078 413 5082 419
rect 5111 413 5114 419
rect 5067 402 5071 409
rect 5037 398 5060 402
rect 5067 399 5082 402
rect 4786 368 4790 397
rect 4811 390 4814 392
rect 4819 390 4822 392
rect 4811 389 4822 390
rect 4804 385 4832 389
rect 4804 379 4808 385
rect 4828 379 4832 385
rect 4817 368 4821 375
rect 4786 364 4810 368
rect 4817 365 4832 368
rect 4828 362 4832 365
rect 4780 356 4821 360
rect 4828 358 4856 362
rect 4828 348 4832 358
rect 4470 345 4724 348
rect 4805 335 4809 344
rect 4805 332 4827 335
rect 4816 331 4827 332
rect 4816 330 4818 331
rect 4822 330 4827 331
rect 4852 289 4856 358
rect 4253 285 4856 289
rect 3434 258 4074 262
rect 1738 254 3223 257
rect 3220 252 3223 254
rect 3220 251 3550 252
rect 3220 249 3554 251
rect 1618 244 2134 247
rect 2131 240 2134 244
rect 2131 238 4328 240
rect 2131 237 4332 238
rect 5037 216 5040 398
rect 5078 396 5082 399
rect 5053 390 5071 394
rect 5078 393 5083 396
rect 5127 393 5130 408
rect 5161 394 5164 740
rect 5182 693 5211 695
rect 5240 695 5243 740
rect 5215 693 5222 695
rect 5182 691 5222 693
rect 5182 667 5186 691
rect 5182 636 5186 663
rect 5191 667 5195 688
rect 5199 684 5214 688
rect 5210 667 5214 684
rect 5191 636 5195 663
rect 5201 636 5205 663
rect 5210 636 5214 663
rect 5218 651 5222 691
rect 5226 681 5233 683
rect 5237 681 5249 683
rect 5226 679 5249 681
rect 5226 667 5230 679
rect 5245 667 5249 679
rect 5218 647 5228 651
rect 5235 643 5239 663
rect 5254 651 5258 663
rect 5246 647 5247 651
rect 5254 647 5257 651
rect 5218 639 5239 643
rect 5201 629 5205 632
rect 5218 629 5222 639
rect 5235 636 5239 639
rect 5254 636 5258 647
rect 5201 625 5222 629
rect 5226 629 5230 632
rect 5245 630 5249 632
rect 5244 629 5249 630
rect 5226 625 5249 629
rect 5226 450 5230 625
rect 5261 529 5291 533
rect 5295 529 5301 533
rect 5261 505 5265 529
rect 5261 474 5265 501
rect 5270 522 5293 526
rect 5270 505 5274 522
rect 5289 505 5293 522
rect 5270 474 5274 501
rect 5280 474 5284 501
rect 5289 474 5293 501
rect 5297 489 5301 529
rect 5305 519 5311 521
rect 5318 521 5321 522
rect 5315 519 5328 521
rect 5305 517 5328 519
rect 5305 505 5309 517
rect 5324 505 5328 517
rect 5297 485 5307 489
rect 5314 481 5318 501
rect 5333 489 5337 501
rect 5325 485 5326 489
rect 5333 485 5336 489
rect 5297 477 5318 481
rect 5280 467 5284 470
rect 5297 467 5301 477
rect 5314 474 5318 477
rect 5333 474 5337 485
rect 5437 478 5449 479
rect 5280 463 5301 467
rect 5427 476 5470 478
rect 5474 477 5520 478
rect 5474 476 5533 477
rect 5427 474 5533 476
rect 5305 467 5309 470
rect 5324 469 5328 470
rect 5321 467 5328 469
rect 5305 466 5328 467
rect 5304 463 5328 466
rect 5427 468 5431 474
rect 5451 468 5455 474
rect 5505 473 5533 474
rect 5505 467 5509 473
rect 5529 467 5533 473
rect 5171 449 5230 450
rect 5318 449 5322 463
rect 5440 457 5444 464
rect 5171 447 5322 449
rect 5171 445 5308 447
rect 5312 445 5322 447
rect 5401 453 5433 457
rect 5440 454 5455 457
rect 5518 456 5522 463
rect 5219 423 5231 424
rect 5209 421 5248 423
rect 5253 421 5269 423
rect 5209 419 5269 421
rect 5273 419 5298 423
rect 5209 413 5213 419
rect 5233 413 5237 419
rect 5266 413 5269 419
rect 5222 402 5226 409
rect 5208 398 5215 402
rect 5222 399 5237 402
rect 5233 396 5237 399
rect 5078 389 5118 393
rect 5127 390 5153 393
rect 5161 390 5226 394
rect 5233 393 5238 396
rect 5282 394 5285 408
rect 5078 382 5082 389
rect 5055 369 5059 378
rect 5127 374 5130 390
rect 5055 368 5087 369
rect 5111 368 5115 369
rect 5055 367 5115 368
rect 5055 366 5094 367
rect 5083 365 5094 366
rect 5098 365 5115 367
rect 5150 342 5153 390
rect 5233 389 5273 393
rect 5282 390 5287 394
rect 5233 382 5237 389
rect 5210 369 5214 378
rect 5282 374 5285 390
rect 5210 367 5239 369
rect 5266 367 5270 369
rect 5210 366 5270 367
rect 5235 364 5245 366
rect 5249 364 5270 366
rect 5401 342 5404 453
rect 5426 449 5429 453
rect 5451 451 5455 454
rect 5503 452 5511 456
rect 5518 453 5533 456
rect 5426 445 5444 449
rect 5451 448 5456 451
rect 5503 448 5507 452
rect 5529 450 5533 453
rect 5529 448 5534 450
rect 5451 444 5463 448
rect 5503 444 5522 448
rect 5529 445 5541 448
rect 5451 437 5455 444
rect 5428 424 5432 433
rect 5428 421 5457 424
rect 5434 419 5435 421
rect 5439 419 5442 421
rect 5460 354 5463 444
rect 5529 436 5533 445
rect 5506 423 5510 432
rect 5506 420 5535 423
rect 5515 418 5517 420
rect 5521 418 5523 420
rect 5538 394 5541 445
rect 5466 391 5541 394
rect 5466 362 5470 391
rect 5491 384 5493 386
rect 5497 384 5502 386
rect 5491 383 5502 384
rect 5484 379 5512 383
rect 5484 373 5488 379
rect 5508 373 5512 379
rect 5497 362 5501 369
rect 5466 358 5490 362
rect 5497 359 5512 362
rect 5508 356 5512 359
rect 5460 350 5501 354
rect 5508 352 5520 356
rect 5508 342 5512 352
rect 5150 339 5404 342
rect 5485 329 5489 338
rect 5485 326 5514 329
rect 5496 324 5501 326
rect 5505 324 5507 326
rect 1502 213 5040 216
rect 1939 202 5174 205
rect 1084 199 1130 202
rect 1112 198 1130 199
rect 1140 198 1144 202
rect 1755 201 5174 202
rect 1112 196 1144 198
rect 1112 194 1124 196
rect 1128 194 1144 196
rect 1410 200 5174 201
rect 1410 198 1944 200
rect 1410 196 1757 198
rect 1410 177 1415 196
rect 1383 173 1415 177
rect 1425 185 1461 187
rect 1465 185 1485 187
rect 1425 183 1485 185
rect 1489 183 1514 187
rect 1425 177 1429 183
rect 1449 177 1453 183
rect 1482 177 1485 183
rect 1081 154 1118 156
rect 1122 154 1141 156
rect 1081 152 1141 154
rect 1145 152 1170 156
rect 1081 146 1085 152
rect 1105 146 1109 152
rect 1138 146 1141 152
rect 1094 135 1098 142
rect 1081 131 1087 135
rect 1094 132 1109 135
rect 1105 129 1109 132
rect 957 114 989 118
rect 998 115 1066 118
rect 1071 123 1098 127
rect 1105 126 1110 129
rect 1154 126 1157 141
rect 1383 126 1387 173
rect 1410 166 1415 173
rect 1438 166 1442 173
rect 1410 162 1431 166
rect 1438 163 1453 166
rect 1424 154 1442 158
rect 1449 157 1453 163
rect 1498 157 1501 172
rect 1520 168 1525 196
rect 1536 187 1572 189
rect 1576 187 1596 189
rect 1536 185 1596 187
rect 1600 185 1625 189
rect 1536 179 1540 185
rect 1560 179 1564 185
rect 1593 179 1596 185
rect 1549 168 1553 175
rect 1520 164 1542 168
rect 1549 165 1564 168
rect 1560 162 1564 165
rect 1449 153 1489 157
rect 1498 153 1509 157
rect 1535 156 1553 160
rect 1560 159 1565 162
rect 1609 159 1612 174
rect 1638 168 1643 196
rect 1652 187 1688 189
rect 1692 187 1712 189
rect 1652 185 1712 187
rect 1716 185 1741 189
rect 1652 179 1656 185
rect 1676 179 1680 185
rect 1709 179 1712 185
rect 1665 168 1669 175
rect 1638 164 1658 168
rect 1665 165 1680 168
rect 1676 162 1680 165
rect 1449 146 1453 153
rect 1426 133 1430 142
rect 1498 138 1501 153
rect 1426 130 1472 133
rect 1482 130 1486 133
rect 1454 129 1486 130
rect 1454 127 1464 129
rect 957 72 961 114
rect 998 99 1001 115
rect 982 87 986 94
rect 972 83 1014 87
rect 972 81 989 83
rect 994 81 1014 83
rect 1071 72 1075 123
rect 1105 122 1145 126
rect 1154 122 1387 126
rect 1468 127 1486 129
rect 1105 115 1109 122
rect 1082 102 1086 111
rect 1154 107 1157 122
rect 1082 100 1128 102
rect 1138 100 1142 102
rect 1082 99 1142 100
rect 1110 97 1128 99
rect 1132 97 1142 99
rect 1366 82 1389 87
rect 957 68 1075 72
rect 1055 38 1059 68
rect 1082 65 1119 67
rect 1123 65 1142 67
rect 1082 63 1142 65
rect 1146 63 1171 67
rect 1082 57 1086 63
rect 1106 57 1110 63
rect 1139 57 1142 63
rect 1095 46 1099 53
rect 1082 42 1088 46
rect 1095 43 1110 46
rect 1106 40 1110 43
rect 1055 34 1099 38
rect 1106 37 1111 40
rect 1106 33 1146 37
rect 1155 34 1158 52
rect 1505 39 1509 153
rect 1560 155 1600 159
rect 1609 156 1618 159
rect 1651 156 1669 160
rect 1676 159 1681 162
rect 1725 159 1728 174
rect 1752 169 1757 196
rect 1772 188 1808 190
rect 1812 188 1832 190
rect 1772 186 1832 188
rect 1836 186 1861 190
rect 1772 180 1776 186
rect 1796 180 1800 186
rect 1829 180 1832 186
rect 1785 169 1789 176
rect 1752 165 1778 169
rect 1785 166 1800 169
rect 1796 163 1800 166
rect 1560 148 1564 155
rect 1537 135 1541 144
rect 1609 140 1612 156
rect 1537 132 1583 135
rect 1593 132 1597 135
rect 1565 131 1597 132
rect 1565 129 1574 131
rect 1578 129 1597 131
rect 1615 45 1618 156
rect 1676 155 1716 159
rect 1725 155 1736 159
rect 1771 157 1789 161
rect 1796 160 1801 163
rect 1845 160 1848 175
rect 1939 170 1944 198
rect 1954 189 1991 191
rect 1995 189 2014 191
rect 1954 187 2014 189
rect 2018 187 2043 191
rect 1954 181 1958 187
rect 1978 181 1982 187
rect 2011 181 2014 187
rect 1967 170 1971 177
rect 1939 166 1960 170
rect 1967 167 1982 170
rect 1676 148 1680 155
rect 1653 135 1657 144
rect 1725 140 1728 155
rect 1653 132 1699 135
rect 1709 132 1713 135
rect 1681 131 1713 132
rect 1681 129 1691 131
rect 1695 129 1713 131
rect 1732 55 1736 155
rect 1796 156 1836 160
rect 1845 156 1880 160
rect 1953 158 1971 162
rect 1978 161 1982 167
rect 2027 161 2030 176
rect 2049 172 2054 200
rect 2065 191 2104 193
rect 2108 191 2125 193
rect 2065 189 2125 191
rect 2129 189 2154 193
rect 2065 183 2069 189
rect 2089 183 2093 189
rect 2122 183 2125 189
rect 2078 172 2082 179
rect 2049 168 2071 172
rect 2078 169 2093 172
rect 2089 166 2093 169
rect 1796 149 1800 156
rect 1773 136 1777 145
rect 1845 141 1848 156
rect 1773 133 1819 136
rect 1829 133 1833 136
rect 1801 132 1833 133
rect 1801 130 1811 132
rect 1815 130 1833 132
rect 1876 63 1880 156
rect 1978 157 2018 161
rect 2027 157 2033 161
rect 2064 160 2082 164
rect 2089 163 2094 166
rect 2138 163 2141 178
rect 2167 172 2172 200
rect 2181 191 2219 193
rect 2223 191 2241 193
rect 2181 189 2241 191
rect 2245 189 2270 193
rect 2181 183 2185 189
rect 2205 183 2209 189
rect 2238 183 2241 189
rect 2194 172 2198 179
rect 2167 168 2187 172
rect 2194 169 2209 172
rect 2205 166 2209 169
rect 2089 159 2129 163
rect 1978 150 1982 157
rect 1955 137 1959 146
rect 2027 142 2030 157
rect 2089 152 2093 159
rect 2138 158 2143 163
rect 2180 160 2198 164
rect 2205 163 2210 166
rect 2254 163 2257 178
rect 2284 173 2289 200
rect 2301 192 2339 194
rect 2343 192 2361 194
rect 2301 190 2361 192
rect 2365 190 2390 194
rect 2301 184 2305 190
rect 2325 184 2329 190
rect 2358 184 2361 190
rect 2314 173 2318 180
rect 2284 169 2307 173
rect 2314 170 2329 173
rect 2325 167 2329 170
rect 2205 159 2245 163
rect 2254 159 2260 163
rect 2300 161 2318 165
rect 2325 164 2330 167
rect 2374 164 2377 179
rect 2325 160 2365 164
rect 2374 160 2380 164
rect 2066 139 2070 148
rect 2138 144 2141 158
rect 2205 152 2209 159
rect 2182 139 2186 148
rect 2254 144 2257 159
rect 2325 153 2329 160
rect 2302 140 2306 149
rect 2374 145 2377 160
rect 1955 134 2001 137
rect 2011 134 2015 137
rect 2066 136 2112 139
rect 2122 136 2126 139
rect 2182 136 2228 139
rect 2238 136 2242 139
rect 2302 137 2348 140
rect 2358 137 2362 140
rect 1983 133 2015 134
rect 2094 135 2126 136
rect 2094 133 2105 135
rect 1983 131 1993 133
rect 1997 131 2015 133
rect 2109 133 2126 135
rect 2210 135 2242 136
rect 2210 133 2220 135
rect 2224 133 2242 135
rect 2330 136 2362 137
rect 2330 134 2341 136
rect 2345 134 2362 136
rect 1876 59 2692 63
rect 1732 51 2676 55
rect 1615 42 2662 45
rect 1505 35 2648 39
rect 1106 26 1110 33
rect 1155 31 1366 34
rect 1083 13 1087 22
rect 1155 18 1158 31
rect 1083 11 1129 13
rect 1139 11 1143 13
rect 1083 10 1143 11
rect 1111 9 1143 10
rect 1363 12 1366 31
rect 1435 21 2311 24
rect 1435 19 1782 21
rect 1435 12 1440 19
rect 1363 9 1440 12
rect 1111 7 1124 9
rect 1128 7 1143 9
rect 1435 -11 1440 9
rect 1450 8 1486 10
rect 1490 8 1510 10
rect 1450 6 1510 8
rect 1514 6 1539 10
rect 1450 2 1454 6
rect 1474 2 1478 6
rect 1507 1 1510 6
rect 1463 -11 1467 -2
rect 1435 -15 1456 -11
rect 1463 -14 1478 -11
rect 1449 -23 1467 -19
rect 1474 -20 1478 -14
rect 1523 -20 1526 -3
rect 1545 -9 1550 19
rect 1561 10 1597 12
rect 1601 10 1621 12
rect 1561 8 1621 10
rect 1625 8 1650 12
rect 1561 2 1565 8
rect 1585 2 1589 8
rect 1618 1 1621 8
rect 1574 -9 1578 -2
rect 1545 -13 1567 -9
rect 1574 -12 1589 -9
rect 1585 -15 1589 -12
rect 1474 -24 1514 -20
rect 1523 -23 1536 -20
rect 1560 -21 1578 -17
rect 1585 -18 1590 -15
rect 1634 -17 1637 -3
rect 1663 -9 1668 19
rect 1677 10 1712 12
rect 1716 10 1737 12
rect 1677 8 1737 10
rect 1741 8 1766 12
rect 1677 2 1681 8
rect 1701 2 1705 8
rect 1734 0 1737 8
rect 1690 -9 1694 -2
rect 1663 -13 1683 -9
rect 1690 -12 1705 -9
rect 1474 -31 1478 -24
rect 1451 -44 1455 -35
rect 1523 -39 1526 -23
rect 833 -49 1124 -47
rect 1451 -47 1497 -44
rect 1507 -47 1511 -44
rect 1128 -49 1228 -47
rect 833 -54 1228 -49
rect 1479 -48 1511 -47
rect 1479 -50 1489 -48
rect 1493 -50 1511 -48
rect 1366 -69 1389 -64
rect 1533 -152 1536 -23
rect 1585 -22 1625 -18
rect 1634 -21 1654 -17
rect 1676 -21 1694 -17
rect 1701 -18 1705 -12
rect 1750 -18 1753 -4
rect 1777 -8 1782 19
rect 1797 11 1834 13
rect 1838 11 1857 13
rect 1797 9 1857 11
rect 1861 9 1886 13
rect 1797 3 1801 9
rect 1821 3 1825 9
rect 1854 0 1857 9
rect 1810 -8 1814 -1
rect 1777 -12 1803 -8
rect 1810 -11 1825 -8
rect 1821 -14 1825 -11
rect 1585 -29 1589 -22
rect 1562 -42 1566 -33
rect 1634 -37 1637 -21
rect 1562 -45 1608 -42
rect 1618 -45 1622 -42
rect 1590 -46 1622 -45
rect 1590 -48 1600 -46
rect 1604 -48 1622 -46
rect 1650 -110 1654 -21
rect 1701 -22 1741 -18
rect 1750 -22 1777 -18
rect 1796 -20 1814 -16
rect 1821 -17 1826 -14
rect 1870 -17 1873 -4
rect 1964 -7 1969 21
rect 1979 12 2016 14
rect 2020 12 2039 14
rect 1979 10 2039 12
rect 2043 10 2068 14
rect 1979 5 1983 10
rect 2003 5 2007 10
rect 2036 4 2039 10
rect 1992 -7 1996 1
rect 1964 -11 1985 -7
rect 1992 -10 2007 -7
rect 1701 -29 1705 -22
rect 1678 -42 1682 -33
rect 1750 -37 1753 -22
rect 1678 -45 1724 -42
rect 1734 -45 1738 -42
rect 1706 -46 1738 -45
rect 1706 -48 1715 -46
rect 1719 -48 1738 -46
rect 1773 -81 1777 -22
rect 1821 -21 1861 -17
rect 1870 -21 1962 -17
rect 1978 -19 1996 -15
rect 2003 -16 2007 -10
rect 2052 -16 2055 0
rect 2074 -5 2079 21
rect 2090 14 2128 16
rect 2132 14 2150 16
rect 2090 12 2150 14
rect 2154 12 2179 16
rect 2090 7 2094 12
rect 2114 7 2118 12
rect 2147 7 2150 12
rect 2103 -5 2107 3
rect 2074 -9 2096 -5
rect 2103 -8 2118 -5
rect 1821 -28 1825 -21
rect 1798 -41 1802 -32
rect 1870 -36 1873 -21
rect 1798 -44 1844 -41
rect 1854 -44 1858 -41
rect 1826 -45 1858 -44
rect 1826 -47 1836 -45
rect 1840 -47 1858 -45
rect 1773 -85 1942 -81
rect 1650 -114 1821 -110
rect 1727 -131 1732 -130
rect 1717 -133 1755 -131
rect 1759 -133 1777 -131
rect 1717 -135 1777 -133
rect 1781 -135 1806 -131
rect 1717 -141 1721 -135
rect 1741 -141 1745 -135
rect 1774 -141 1777 -135
rect 1730 -152 1734 -145
rect 1533 -156 1723 -152
rect 1730 -155 1745 -152
rect 1741 -158 1745 -155
rect 1716 -164 1734 -160
rect 1741 -161 1746 -158
rect 1790 -161 1793 -146
rect 1817 -153 1821 -114
rect 1845 -132 1850 -131
rect 1835 -134 1871 -132
rect 1875 -134 1895 -132
rect 1835 -136 1895 -134
rect 1899 -136 1924 -132
rect 1835 -142 1839 -136
rect 1859 -142 1863 -136
rect 1892 -142 1895 -136
rect 1848 -153 1852 -146
rect 1817 -157 1841 -153
rect 1848 -156 1863 -153
rect 1859 -159 1863 -156
rect 1741 -165 1781 -161
rect 1790 -164 1795 -161
rect 1741 -172 1745 -165
rect 1718 -185 1722 -176
rect 1790 -180 1793 -164
rect 1823 -165 1852 -161
rect 1859 -162 1864 -159
rect 1908 -162 1911 -147
rect 1938 -153 1942 -85
rect 1958 -120 1962 -21
rect 2003 -20 2043 -16
rect 2052 -20 2066 -16
rect 2089 -17 2107 -13
rect 2114 -14 2118 -8
rect 2163 -14 2166 3
rect 2192 -5 2197 21
rect 2206 14 2245 16
rect 2249 14 2266 16
rect 2206 12 2266 14
rect 2270 12 2295 16
rect 2206 7 2210 12
rect 2230 7 2234 12
rect 2263 6 2266 12
rect 2219 -5 2223 3
rect 2192 -9 2212 -5
rect 2219 -8 2234 -5
rect 2003 -27 2007 -20
rect 1980 -40 1984 -31
rect 2052 -35 2055 -20
rect 1980 -43 2026 -40
rect 2036 -43 2040 -40
rect 2008 -44 2040 -43
rect 2008 -46 2018 -44
rect 2022 -46 2040 -44
rect 2062 -61 2066 -20
rect 2114 -18 2154 -14
rect 2163 -18 2186 -14
rect 2205 -17 2223 -13
rect 2230 -14 2234 -8
rect 2279 -14 2282 3
rect 2306 -5 2311 21
rect 2326 15 2364 17
rect 2368 15 2386 17
rect 2326 13 2386 15
rect 2390 13 2415 17
rect 2326 7 2330 13
rect 2350 7 2354 13
rect 2383 7 2386 13
rect 2339 -4 2343 3
rect 2306 -8 2332 -5
rect 2339 -7 2354 -4
rect 2114 -25 2118 -18
rect 2091 -38 2095 -29
rect 2163 -33 2166 -18
rect 2091 -41 2137 -38
rect 2147 -41 2151 -38
rect 2119 -42 2151 -41
rect 2119 -44 2129 -42
rect 2133 -44 2151 -42
rect 2182 -50 2186 -18
rect 2230 -18 2270 -14
rect 2279 -17 2290 -14
rect 2327 -16 2343 -12
rect 2350 -13 2354 -7
rect 2399 -13 2402 3
rect 2230 -25 2234 -18
rect 2207 -38 2211 -29
rect 2279 -33 2282 -17
rect 2207 -41 2253 -38
rect 2263 -41 2267 -38
rect 2235 -42 2267 -41
rect 2235 -44 2245 -42
rect 2249 -44 2267 -42
rect 1958 -124 2072 -120
rect 1978 -132 1983 -131
rect 1968 -135 2004 -132
rect 2009 -135 2028 -132
rect 1968 -136 2028 -135
rect 2032 -136 2057 -132
rect 1968 -142 1972 -136
rect 1992 -142 1996 -136
rect 2025 -142 2028 -136
rect 1981 -153 1985 -146
rect 1938 -157 1974 -153
rect 1981 -156 1996 -153
rect 1992 -159 1996 -156
rect 1859 -166 1899 -162
rect 1908 -165 1913 -162
rect 1967 -165 1985 -161
rect 1992 -162 1997 -159
rect 2041 -162 2044 -147
rect 2068 -154 2072 -124
rect 2097 -133 2102 -132
rect 2087 -135 2124 -133
rect 2128 -135 2147 -133
rect 2087 -137 2147 -135
rect 2151 -137 2176 -133
rect 2087 -143 2091 -137
rect 2111 -143 2115 -137
rect 2144 -143 2147 -137
rect 2100 -154 2104 -147
rect 2068 -158 2093 -154
rect 2100 -157 2115 -154
rect 2111 -160 2115 -157
rect 1859 -173 1863 -166
rect 1718 -187 1764 -185
rect 1774 -187 1778 -185
rect 1718 -188 1778 -187
rect 1746 -190 1754 -188
rect 1758 -190 1778 -188
rect 1836 -186 1840 -177
rect 1908 -181 1911 -165
rect 1992 -166 2032 -162
rect 2041 -165 2046 -162
rect 1992 -173 1996 -166
rect 1969 -186 1973 -177
rect 2041 -181 2044 -165
rect 2073 -166 2104 -162
rect 2111 -163 2116 -160
rect 2160 -163 2163 -148
rect 1836 -189 1882 -186
rect 1864 -190 1882 -189
rect 1892 -190 1896 -186
rect 1969 -189 2015 -186
rect 1864 -192 1896 -190
rect 1864 -194 1873 -192
rect 1877 -194 1896 -192
rect 1997 -190 2015 -189
rect 2025 -190 2029 -186
rect 1997 -191 2029 -190
rect 1997 -193 2006 -191
rect 2010 -193 2029 -191
rect 2073 -216 2077 -166
rect 2111 -167 2151 -163
rect 2160 -166 2165 -163
rect 2111 -174 2115 -167
rect 2088 -187 2092 -178
rect 2160 -182 2163 -166
rect 2088 -190 2134 -187
rect 2144 -190 2148 -187
rect 2116 -191 2148 -190
rect 2116 -193 2122 -191
rect 2126 -193 2148 -191
rect 2287 -204 2290 -17
rect 2350 -17 2390 -13
rect 2399 -17 2435 -13
rect 2350 -24 2354 -17
rect 2327 -37 2331 -28
rect 2399 -32 2402 -17
rect 2327 -40 2373 -37
rect 2383 -40 2387 -37
rect 2355 -41 2387 -40
rect 2355 -43 2366 -41
rect 2370 -43 2387 -41
rect 2431 -216 2435 -17
rect 2073 -220 2435 -216
rect 2644 -611 2648 35
rect 2659 -568 2662 42
rect 2672 -551 2676 51
rect 2688 -530 2692 59
rect 3595 26 3600 27
rect 3585 24 3631 26
rect 3635 25 3678 26
rect 3635 24 3691 25
rect 3585 22 3691 24
rect 3585 16 3589 22
rect 3609 16 3613 22
rect 3663 21 3691 22
rect 3663 15 3667 21
rect 3687 15 3691 21
rect 3598 5 3602 12
rect 3581 1 3591 5
rect 3598 2 3613 5
rect 3676 4 3680 11
rect 3584 -3 3587 1
rect 3584 -7 3592 -3
rect 3595 -7 3602 -3
rect 3609 -5 3613 2
rect 3661 0 3669 4
rect 3676 0 3691 4
rect 3661 -1 3670 0
rect 3663 -5 3666 -1
rect 3687 -4 3691 0
rect 3609 -8 3621 -5
rect 3663 -8 3680 -5
rect 3687 -7 3699 -4
rect 3609 -15 3613 -8
rect 3586 -28 3590 -19
rect 3586 -31 3615 -28
rect 3595 -33 3602 -31
rect 3618 -98 3621 -8
rect 3687 -16 3691 -7
rect 3664 -29 3668 -20
rect 3664 -31 3693 -29
rect 3664 -32 3681 -31
rect 3675 -34 3681 -32
rect 3685 -32 3693 -31
rect 3696 -58 3699 -7
rect 3624 -61 3699 -58
rect 3624 -90 3628 -61
rect 3652 -68 3654 -66
rect 3658 -68 3659 -66
rect 3652 -69 3659 -68
rect 3642 -73 3670 -69
rect 3642 -79 3646 -73
rect 3666 -79 3670 -73
rect 3655 -90 3659 -83
rect 3624 -94 3648 -90
rect 3655 -93 3670 -90
rect 3666 -96 3670 -93
rect 3618 -102 3659 -98
rect 3666 -100 3672 -96
rect 3666 -110 3670 -100
rect 3813 -101 3818 -100
rect 3803 -103 3839 -101
rect 3843 -102 3896 -101
rect 3843 -103 3909 -102
rect 3803 -105 3909 -103
rect 3803 -111 3807 -105
rect 3827 -111 3831 -105
rect 3643 -123 3647 -114
rect 3881 -106 3909 -105
rect 3881 -112 3885 -106
rect 3905 -112 3909 -106
rect 3816 -122 3820 -115
rect 3643 -126 3672 -123
rect 3779 -126 3809 -122
rect 3816 -125 3831 -122
rect 3894 -123 3898 -116
rect 3654 -127 3662 -126
rect 3654 -128 3656 -127
rect 3660 -128 3662 -127
rect 2786 -215 2827 -211
rect 3608 -250 3613 -249
rect 3598 -252 3649 -250
rect 3653 -251 3691 -250
rect 3653 -252 3704 -251
rect 3598 -254 3704 -252
rect 3598 -260 3602 -254
rect 3622 -260 3626 -254
rect 3676 -255 3704 -254
rect 3676 -261 3680 -255
rect 3700 -261 3704 -255
rect 3611 -271 3615 -264
rect 3594 -275 3604 -271
rect 3611 -274 3626 -271
rect 3689 -272 3693 -265
rect 3597 -279 3600 -275
rect 3622 -277 3626 -274
rect 3674 -276 3682 -272
rect 3689 -275 3704 -272
rect 3597 -283 3615 -279
rect 3622 -280 3627 -277
rect 3674 -280 3678 -276
rect 3700 -278 3704 -275
rect 3700 -280 3705 -278
rect 3622 -284 3634 -280
rect 3674 -284 3693 -280
rect 3700 -283 3712 -280
rect 3622 -291 3626 -284
rect 3599 -304 3603 -295
rect 3599 -307 3628 -304
rect 3608 -309 3610 -307
rect 3614 -309 3615 -307
rect 3631 -374 3634 -284
rect 3700 -292 3704 -283
rect 3677 -305 3681 -296
rect 3677 -307 3706 -305
rect 3677 -308 3694 -307
rect 3688 -310 3694 -308
rect 3698 -308 3706 -307
rect 3709 -334 3712 -283
rect 3637 -337 3712 -334
rect 3637 -366 3641 -337
rect 3665 -344 3666 -342
rect 3670 -344 3672 -342
rect 3665 -345 3674 -344
rect 3655 -349 3683 -345
rect 3655 -355 3659 -349
rect 3679 -355 3683 -349
rect 3668 -366 3672 -359
rect 3637 -370 3661 -366
rect 3668 -369 3683 -366
rect 3679 -372 3683 -369
rect 3779 -372 3783 -126
rect 3802 -130 3805 -126
rect 3827 -128 3831 -125
rect 3879 -127 3887 -123
rect 3894 -126 3909 -123
rect 3802 -134 3820 -130
rect 3827 -131 3832 -128
rect 3879 -131 3883 -127
rect 3905 -129 3909 -126
rect 3905 -131 3910 -129
rect 3827 -135 3839 -131
rect 3879 -135 3898 -131
rect 3905 -134 3917 -131
rect 3827 -142 3831 -135
rect 3804 -155 3808 -146
rect 3804 -158 3833 -155
rect 3813 -160 3815 -158
rect 3819 -160 3820 -158
rect 3836 -225 3839 -135
rect 3905 -143 3909 -134
rect 3882 -156 3886 -147
rect 3882 -158 3911 -156
rect 3882 -159 3904 -158
rect 3893 -161 3899 -159
rect 3908 -159 3911 -158
rect 3914 -185 3917 -134
rect 4086 -142 4099 -138
rect 4103 -140 4108 -138
rect 4112 -140 4127 -138
rect 4103 -142 4127 -140
rect 4096 -148 4099 -142
rect 4112 -168 4115 -153
rect 3842 -188 3917 -185
rect 3998 -172 4103 -168
rect 4112 -171 4901 -168
rect 3842 -217 3846 -188
rect 3870 -195 3871 -193
rect 3875 -195 3877 -193
rect 3870 -196 3877 -195
rect 3860 -200 3888 -196
rect 3860 -206 3864 -200
rect 3884 -206 3888 -200
rect 3873 -217 3877 -210
rect 3842 -221 3866 -217
rect 3873 -220 3888 -217
rect 3884 -223 3888 -220
rect 3998 -223 4002 -172
rect 4112 -187 4115 -171
rect 4096 -199 4100 -192
rect 4086 -203 4128 -199
rect 4086 -205 4106 -203
rect 4110 -205 4128 -203
rect 3836 -229 3877 -225
rect 3884 -227 4002 -223
rect 3884 -237 3888 -227
rect 3861 -250 3865 -241
rect 3861 -253 3890 -250
rect 3872 -255 3874 -253
rect 3878 -255 3880 -253
rect 3631 -378 3672 -374
rect 3679 -376 3783 -372
rect 3679 -386 3683 -376
rect 3656 -399 3660 -390
rect 3656 -402 3685 -399
rect 3667 -404 3669 -402
rect 3673 -404 3675 -402
rect 2813 -521 4726 -518
rect 2688 -534 2762 -530
rect 2672 -555 2764 -551
rect 2659 -571 2764 -568
rect 2644 -616 2764 -611
rect 2712 -669 2806 -665
rect 2713 -682 2792 -678
rect 2715 -696 2773 -692
rect 2717 -735 2758 -731
rect 2752 -1243 2756 -735
rect 2765 -1202 2769 -696
rect 2781 -1180 2785 -682
rect 2799 -1165 2803 -669
rect 2813 -868 2816 -521
rect 3656 -578 4136 -576
rect 2819 -586 2832 -582
rect 2836 -584 2841 -582
rect 2845 -584 2860 -582
rect 2836 -586 2860 -584
rect 2984 -586 2997 -582
rect 3001 -584 3004 -582
rect 3008 -584 3025 -582
rect 3001 -586 3025 -584
rect 3161 -585 3174 -581
rect 3178 -583 3183 -581
rect 3656 -580 4132 -578
rect 3187 -583 3202 -581
rect 3178 -585 3202 -583
rect 2829 -592 2832 -586
rect 2994 -592 2997 -586
rect 3171 -591 3174 -585
rect 3336 -586 3349 -582
rect 3353 -584 3358 -582
rect 3362 -584 3377 -582
rect 3353 -586 3377 -584
rect 2845 -612 2848 -597
rect 3010 -612 3013 -597
rect 3187 -611 3190 -596
rect 3346 -592 3349 -586
rect 2835 -616 2836 -612
rect 2845 -615 2866 -612
rect 2845 -631 2848 -615
rect 2829 -643 2833 -636
rect 2825 -648 2856 -643
rect 2825 -649 2834 -648
rect 2838 -649 2856 -648
rect 2842 -817 2846 -736
rect 2850 -764 2856 -649
rect 2863 -722 2866 -615
rect 3000 -616 3001 -612
rect 3010 -615 3037 -612
rect 3176 -615 3178 -611
rect 3187 -614 3230 -611
rect 3362 -612 3365 -597
rect 3010 -631 3013 -615
rect 2994 -643 2998 -636
rect 2984 -648 3026 -643
rect 2984 -649 3001 -648
rect 3006 -649 3026 -648
rect 2885 -701 2890 -700
rect 2875 -703 2911 -701
rect 2915 -703 2935 -701
rect 2875 -705 2935 -703
rect 2939 -705 2964 -701
rect 2875 -711 2879 -705
rect 2899 -711 2903 -705
rect 2932 -711 2935 -705
rect 2888 -722 2892 -715
rect 2863 -726 2881 -722
rect 2888 -725 2903 -722
rect 2899 -728 2903 -725
rect 2874 -734 2892 -730
rect 2899 -731 2904 -728
rect 2948 -731 2951 -716
rect 3034 -717 3037 -615
rect 3187 -630 3190 -614
rect 3171 -642 3175 -635
rect 3161 -647 3203 -642
rect 3161 -648 3178 -647
rect 3183 -648 3203 -647
rect 3056 -696 3061 -695
rect 3046 -698 3085 -696
rect 3089 -698 3106 -696
rect 3046 -700 3106 -698
rect 3110 -700 3135 -696
rect 3046 -706 3050 -700
rect 3070 -706 3074 -700
rect 3103 -706 3106 -700
rect 3059 -717 3063 -710
rect 3034 -721 3052 -717
rect 3059 -720 3074 -717
rect 3070 -723 3074 -720
rect 3045 -729 3063 -725
rect 3070 -726 3075 -723
rect 3119 -725 3122 -711
rect 3227 -721 3230 -614
rect 3352 -616 3353 -612
rect 3362 -615 3411 -612
rect 3362 -631 3365 -615
rect 3346 -643 3350 -636
rect 3341 -648 3378 -643
rect 3341 -649 3353 -648
rect 3357 -649 3378 -648
rect 3249 -700 3254 -699
rect 3239 -702 3275 -700
rect 3279 -702 3299 -700
rect 3239 -704 3299 -702
rect 3303 -704 3328 -700
rect 3239 -710 3243 -704
rect 3263 -710 3267 -704
rect 3296 -710 3299 -704
rect 3252 -721 3256 -714
rect 3227 -725 3245 -721
rect 3252 -724 3267 -721
rect 2899 -735 2939 -731
rect 2948 -734 2967 -731
rect 2899 -742 2903 -735
rect 2876 -755 2880 -746
rect 2948 -750 2951 -734
rect 2876 -758 2922 -755
rect 2932 -758 2936 -755
rect 2879 -764 2885 -758
rect 2904 -760 2936 -758
rect 2904 -761 2913 -760
rect 2917 -761 2936 -760
rect 2850 -770 2885 -764
rect 2842 -821 2956 -817
rect 2964 -861 2967 -734
rect 3021 -792 3025 -731
rect 3070 -730 3110 -726
rect 3119 -729 3123 -725
rect 3263 -727 3267 -724
rect 3070 -737 3074 -730
rect 3047 -750 3051 -741
rect 3119 -745 3122 -729
rect 3239 -733 3256 -729
rect 3263 -730 3268 -727
rect 3312 -730 3315 -715
rect 3408 -717 3411 -615
rect 3430 -696 3435 -695
rect 3420 -698 3457 -696
rect 3461 -698 3480 -696
rect 3420 -700 3480 -698
rect 3484 -700 3509 -696
rect 3420 -706 3424 -700
rect 3444 -706 3448 -700
rect 3477 -706 3480 -700
rect 3433 -717 3437 -710
rect 3408 -721 3426 -717
rect 3433 -720 3448 -717
rect 3444 -723 3448 -720
rect 3419 -729 3437 -725
rect 3444 -726 3449 -723
rect 3493 -725 3496 -711
rect 3444 -730 3484 -726
rect 3493 -729 3497 -725
rect 3047 -753 3093 -750
rect 3103 -753 3107 -750
rect 3075 -755 3107 -753
rect 3075 -756 3085 -755
rect 3089 -756 3107 -755
rect 3210 -782 3214 -735
rect 3263 -734 3303 -730
rect 3312 -734 3324 -730
rect 3263 -741 3267 -734
rect 3240 -754 3244 -745
rect 3312 -749 3315 -734
rect 3444 -737 3448 -730
rect 3421 -750 3425 -741
rect 3493 -745 3496 -729
rect 3421 -753 3467 -750
rect 3477 -753 3481 -750
rect 3240 -757 3286 -754
rect 3296 -757 3300 -754
rect 3449 -755 3481 -753
rect 3449 -756 3458 -755
rect 3268 -759 3300 -757
rect 3462 -756 3481 -755
rect 3268 -760 3277 -759
rect 3281 -760 3300 -759
rect 3656 -782 3660 -580
rect 3210 -786 3660 -782
rect 3682 -588 4379 -587
rect 3682 -591 4375 -588
rect 3682 -792 3686 -591
rect 4462 -591 4649 -589
rect 4462 -593 4645 -591
rect 4462 -596 4466 -593
rect 3021 -796 3686 -792
rect 3701 -600 4466 -596
rect 3701 -817 3705 -600
rect 3734 -631 3747 -627
rect 3751 -629 3754 -627
rect 3826 -626 3862 -623
rect 4225 -623 4238 -619
rect 4242 -621 4247 -619
rect 4317 -619 4346 -615
rect 4350 -619 4357 -615
rect 4494 -618 4507 -614
rect 4511 -616 4514 -614
rect 4586 -613 4618 -610
rect 4622 -613 4626 -610
rect 4586 -614 4626 -613
rect 4518 -616 4535 -614
rect 4511 -618 4535 -616
rect 4251 -621 4266 -619
rect 4242 -623 4266 -621
rect 3826 -627 3866 -626
rect 3758 -629 3775 -627
rect 3751 -631 3775 -629
rect 3744 -637 3747 -631
rect 3760 -656 3763 -642
rect 3826 -651 3830 -627
rect 3750 -661 3751 -657
rect 3760 -659 3793 -656
rect 3760 -676 3763 -659
rect 3744 -688 3748 -681
rect 3734 -692 3776 -688
rect 3734 -694 3737 -692
rect 3741 -693 3776 -692
rect 3741 -694 3751 -693
rect 3756 -694 3776 -693
rect 2988 -821 3705 -817
rect 3790 -789 3793 -659
rect 3826 -682 3830 -655
rect 3835 -634 3838 -630
rect 3842 -634 3858 -630
rect 3835 -651 3839 -634
rect 3854 -651 3858 -634
rect 3835 -682 3839 -655
rect 3845 -682 3849 -655
rect 3854 -682 3858 -655
rect 3862 -667 3866 -627
rect 3982 -632 3995 -628
rect 3999 -630 4003 -628
rect 4074 -627 4105 -624
rect 4109 -627 4114 -624
rect 4074 -628 4114 -627
rect 4007 -630 4023 -628
rect 3999 -632 4023 -630
rect 3870 -637 3878 -635
rect 3883 -637 3893 -635
rect 3870 -639 3893 -637
rect 3870 -651 3874 -639
rect 3889 -651 3893 -639
rect 3992 -638 3995 -632
rect 3862 -671 3872 -667
rect 3879 -675 3883 -655
rect 3898 -667 3902 -655
rect 4008 -658 4011 -643
rect 4074 -652 4078 -628
rect 3998 -662 3999 -658
rect 4008 -662 4010 -658
rect 3890 -672 3891 -668
rect 3898 -671 3901 -667
rect 3862 -679 3883 -675
rect 3845 -689 3849 -686
rect 3862 -689 3866 -679
rect 3879 -682 3883 -679
rect 3898 -682 3902 -671
rect 4008 -677 4011 -662
rect 3845 -693 3866 -689
rect 3870 -689 3874 -686
rect 3889 -689 3893 -686
rect 3992 -689 3996 -682
rect 4074 -683 4078 -656
rect 4083 -635 4086 -631
rect 4090 -635 4106 -631
rect 4083 -652 4087 -635
rect 4102 -652 4106 -635
rect 4083 -683 4087 -656
rect 4093 -683 4097 -656
rect 4102 -683 4106 -656
rect 4110 -668 4114 -628
rect 4235 -629 4238 -623
rect 4118 -638 4125 -636
rect 4129 -638 4141 -636
rect 4118 -640 4141 -638
rect 4118 -652 4122 -640
rect 4137 -652 4141 -640
rect 4241 -653 4242 -649
rect 4251 -650 4254 -634
rect 4317 -643 4321 -619
rect 4251 -653 4294 -650
rect 4110 -672 4120 -668
rect 4127 -676 4131 -656
rect 4146 -668 4150 -656
rect 4251 -668 4254 -653
rect 4138 -672 4139 -668
rect 4146 -672 4149 -668
rect 4110 -680 4131 -676
rect 3870 -693 3875 -689
rect 3879 -690 3893 -689
rect 3982 -690 4024 -689
rect 3879 -693 4024 -690
rect 3983 -695 4024 -693
rect 4093 -690 4097 -687
rect 4110 -690 4114 -680
rect 4127 -683 4131 -680
rect 4146 -683 4150 -672
rect 4235 -680 4239 -673
rect 4093 -694 4114 -690
rect 4217 -685 4267 -680
rect 4217 -686 4244 -685
rect 4118 -690 4122 -687
rect 4137 -690 4141 -687
rect 4118 -694 4141 -690
rect 4006 -702 4012 -695
rect 4123 -702 4129 -694
rect 4217 -702 4223 -686
rect 4248 -686 4267 -685
rect 4006 -706 4223 -702
rect 4010 -708 4223 -706
rect 4291 -748 4294 -653
rect 4317 -674 4321 -647
rect 4326 -626 4329 -622
rect 4333 -626 4349 -622
rect 4326 -643 4330 -626
rect 4345 -643 4349 -626
rect 4326 -674 4330 -647
rect 4336 -674 4340 -647
rect 4345 -674 4349 -647
rect 4353 -659 4357 -619
rect 4504 -624 4507 -618
rect 4361 -629 4363 -627
rect 4367 -629 4384 -627
rect 4361 -631 4384 -629
rect 4361 -643 4365 -631
rect 4380 -643 4384 -631
rect 4353 -663 4363 -659
rect 4370 -667 4374 -647
rect 4389 -659 4393 -647
rect 4510 -648 4511 -644
rect 4381 -663 4382 -659
rect 4389 -663 4392 -659
rect 4520 -663 4523 -629
rect 4353 -671 4374 -667
rect 4336 -681 4340 -678
rect 4353 -681 4357 -671
rect 4370 -674 4374 -671
rect 4389 -674 4393 -663
rect 4336 -685 4357 -681
rect 4586 -638 4590 -614
rect 4504 -675 4508 -668
rect 4586 -669 4590 -642
rect 4595 -621 4598 -617
rect 4602 -621 4618 -617
rect 4595 -638 4599 -621
rect 4614 -638 4618 -621
rect 4595 -669 4599 -642
rect 4605 -669 4609 -642
rect 4614 -669 4618 -642
rect 4622 -654 4626 -614
rect 4630 -624 4634 -622
rect 4638 -624 4653 -622
rect 4630 -626 4653 -624
rect 4630 -638 4634 -626
rect 4649 -638 4653 -626
rect 4622 -658 4632 -654
rect 4639 -662 4643 -642
rect 4658 -654 4662 -642
rect 4650 -658 4651 -654
rect 4658 -658 4661 -654
rect 4622 -666 4643 -662
rect 4504 -678 4536 -675
rect 4361 -681 4365 -678
rect 4380 -681 4384 -678
rect 4510 -681 4536 -678
rect 4605 -676 4609 -673
rect 4622 -676 4626 -666
rect 4639 -669 4643 -666
rect 4658 -669 4662 -658
rect 4605 -680 4626 -676
rect 4630 -676 4634 -673
rect 4649 -676 4653 -673
rect 4630 -680 4653 -676
rect 4361 -685 4369 -681
rect 4373 -685 4516 -681
rect 4512 -690 4516 -685
rect 4639 -690 4643 -680
rect 4512 -694 4643 -690
rect 4291 -751 4437 -748
rect 4088 -757 4093 -756
rect 4078 -759 4115 -757
rect 4119 -759 4138 -757
rect 4078 -761 4138 -759
rect 4142 -761 4167 -757
rect 4078 -767 4082 -761
rect 4102 -767 4106 -761
rect 4135 -767 4138 -761
rect 4091 -778 4095 -771
rect 4074 -782 4084 -779
rect 4091 -781 4106 -778
rect 4102 -784 4106 -781
rect 4085 -787 4095 -786
rect 4062 -789 4095 -787
rect 3790 -790 4095 -789
rect 4102 -787 4107 -784
rect 4151 -787 4154 -772
rect 4242 -769 4427 -766
rect 4242 -787 4245 -769
rect 4308 -777 4313 -776
rect 4298 -779 4335 -777
rect 4339 -779 4358 -777
rect 4298 -781 4358 -779
rect 4362 -781 4387 -777
rect 4298 -787 4302 -781
rect 4322 -787 4326 -781
rect 3790 -792 4068 -790
rect 4102 -791 4142 -787
rect 4151 -790 4251 -787
rect 3017 -840 3022 -839
rect 3007 -842 3045 -840
rect 3049 -842 3067 -840
rect 3007 -844 3067 -842
rect 3071 -844 3096 -840
rect 3007 -850 3011 -844
rect 3031 -850 3035 -844
rect 3064 -850 3067 -844
rect 3020 -861 3024 -854
rect 2964 -865 3013 -861
rect 3020 -864 3035 -861
rect 3031 -867 3035 -864
rect 2813 -869 3015 -868
rect 2813 -873 3024 -869
rect 3031 -870 3036 -867
rect 3080 -869 3083 -855
rect 2977 -1060 2982 -873
rect 3031 -874 3071 -870
rect 3080 -873 3085 -869
rect 3031 -881 3035 -874
rect 3008 -894 3012 -885
rect 3080 -889 3083 -873
rect 3008 -897 3054 -894
rect 3064 -897 3068 -894
rect 3036 -898 3068 -897
rect 3036 -900 3047 -898
rect 3051 -900 3068 -898
rect 3790 -902 3793 -792
rect 4102 -798 4106 -791
rect 4079 -811 4083 -802
rect 4151 -806 4154 -790
rect 4079 -814 4125 -811
rect 4135 -814 4139 -811
rect 4107 -815 4139 -814
rect 4107 -817 4116 -815
rect 4120 -817 4139 -815
rect 3867 -872 3872 -871
rect 3857 -874 3895 -872
rect 3899 -874 3917 -872
rect 3857 -876 3917 -874
rect 3921 -876 3946 -872
rect 3857 -882 3861 -876
rect 3881 -882 3885 -876
rect 3914 -882 3917 -876
rect 3870 -893 3874 -886
rect 3853 -897 3863 -894
rect 3870 -896 3885 -893
rect 3881 -899 3885 -896
rect 3864 -902 3874 -901
rect 3790 -905 3874 -902
rect 3881 -902 3886 -899
rect 3930 -901 3933 -887
rect 3021 -1038 3026 -1037
rect 3011 -1040 3048 -1038
rect 3052 -1040 3071 -1038
rect 3011 -1042 3071 -1040
rect 3075 -1042 3100 -1038
rect 3011 -1048 3015 -1042
rect 3035 -1048 3039 -1042
rect 3068 -1048 3071 -1042
rect 3024 -1059 3028 -1052
rect 2977 -1063 3017 -1060
rect 3024 -1062 3039 -1059
rect 3035 -1065 3039 -1062
rect 3018 -1068 3028 -1067
rect 2995 -1071 3028 -1068
rect 3035 -1068 3040 -1065
rect 3084 -1067 3087 -1053
rect 2799 -1169 2978 -1165
rect 2781 -1184 2978 -1180
rect 2765 -1206 2984 -1202
rect 2844 -1217 2857 -1213
rect 2861 -1215 2864 -1213
rect 2868 -1215 2885 -1213
rect 2861 -1217 2885 -1215
rect 2854 -1223 2857 -1217
rect 2870 -1243 2873 -1228
rect 2980 -1243 2984 -1206
rect 2752 -1247 2861 -1243
rect 2870 -1246 2891 -1243
rect 2870 -1262 2873 -1246
rect 2854 -1274 2858 -1267
rect 2844 -1278 2881 -1274
rect 2844 -1280 2858 -1278
rect 2862 -1280 2881 -1278
rect 2875 -1386 2881 -1280
rect 2888 -1353 2891 -1246
rect 2980 -1247 2982 -1243
rect 2910 -1332 2915 -1331
rect 2900 -1334 2936 -1332
rect 2940 -1334 2960 -1332
rect 2900 -1336 2960 -1334
rect 2964 -1336 2989 -1332
rect 2900 -1342 2904 -1336
rect 2924 -1342 2928 -1336
rect 2957 -1342 2960 -1336
rect 2913 -1353 2917 -1346
rect 2888 -1357 2906 -1353
rect 2913 -1356 2928 -1353
rect 2924 -1359 2928 -1356
rect 2900 -1365 2917 -1361
rect 2924 -1362 2929 -1359
rect 2973 -1362 2976 -1347
rect 2995 -1362 2998 -1071
rect 3035 -1072 3075 -1068
rect 3084 -1071 3089 -1067
rect 3035 -1079 3039 -1072
rect 3012 -1092 3016 -1083
rect 3084 -1087 3087 -1071
rect 3790 -1080 3793 -905
rect 3881 -906 3921 -902
rect 3930 -905 3934 -901
rect 3881 -913 3885 -906
rect 3858 -926 3862 -917
rect 3930 -921 3933 -905
rect 3858 -929 3904 -926
rect 3914 -929 3918 -926
rect 3886 -931 3918 -929
rect 3886 -932 3895 -931
rect 3899 -932 3918 -931
rect 4006 -1026 4010 -1008
rect 3880 -1058 3885 -1057
rect 3870 -1060 3905 -1058
rect 3909 -1060 3930 -1058
rect 3870 -1062 3930 -1060
rect 3934 -1062 3959 -1058
rect 3870 -1068 3874 -1062
rect 3894 -1068 3898 -1062
rect 3927 -1068 3930 -1062
rect 4170 -1063 4173 -790
rect 4248 -807 4251 -790
rect 4355 -787 4358 -781
rect 4311 -798 4315 -791
rect 4294 -802 4304 -799
rect 4311 -801 4326 -798
rect 4322 -804 4326 -801
rect 4305 -807 4315 -806
rect 4248 -810 4315 -807
rect 4322 -807 4327 -804
rect 4371 -806 4374 -792
rect 4424 -799 4427 -769
rect 4434 -791 4437 -751
rect 4464 -769 4469 -768
rect 4454 -771 4489 -769
rect 4493 -771 4514 -769
rect 4454 -773 4514 -771
rect 4518 -773 4543 -769
rect 4454 -779 4458 -773
rect 4478 -779 4482 -773
rect 4511 -779 4514 -773
rect 4467 -790 4471 -783
rect 4434 -794 4460 -791
rect 4467 -793 4482 -790
rect 4478 -796 4482 -793
rect 4461 -799 4471 -798
rect 4424 -802 4471 -799
rect 4478 -799 4483 -796
rect 4527 -799 4530 -784
rect 4723 -799 4726 -521
rect 4478 -803 4518 -799
rect 4527 -802 4726 -799
rect 4322 -811 4362 -807
rect 4371 -810 4376 -806
rect 4478 -810 4482 -803
rect 4322 -818 4326 -811
rect 4299 -831 4303 -822
rect 4371 -826 4374 -810
rect 4455 -823 4459 -814
rect 4527 -818 4530 -802
rect 4455 -826 4501 -823
rect 4511 -826 4515 -823
rect 4483 -827 4515 -826
rect 4483 -829 4492 -827
rect 4496 -829 4515 -827
rect 4299 -834 4345 -831
rect 4355 -834 4359 -831
rect 4327 -835 4359 -834
rect 4327 -837 4336 -835
rect 4340 -837 4359 -835
rect 4898 -1016 4901 -171
rect 5018 -994 5023 -993
rect 5008 -996 5045 -994
rect 5049 -996 5068 -994
rect 5008 -998 5068 -996
rect 5072 -998 5097 -994
rect 5008 -1004 5012 -998
rect 5032 -1004 5036 -998
rect 5065 -1004 5068 -998
rect 5021 -1015 5025 -1008
rect 4898 -1019 5014 -1016
rect 5021 -1018 5036 -1015
rect 5032 -1021 5036 -1018
rect 5015 -1024 5025 -1023
rect 4897 -1027 5025 -1024
rect 5032 -1024 5037 -1021
rect 5081 -1024 5084 -1009
rect 5169 -1017 5174 200
rect 5235 -995 5240 -994
rect 5225 -997 5260 -995
rect 5264 -997 5285 -995
rect 5225 -999 5285 -997
rect 5289 -999 5314 -995
rect 5225 -1005 5229 -999
rect 5249 -1005 5253 -999
rect 5282 -1005 5285 -999
rect 5238 -1016 5242 -1009
rect 5169 -1020 5231 -1017
rect 5238 -1019 5253 -1016
rect 5249 -1022 5253 -1019
rect 4208 -1041 4213 -1040
rect 4198 -1043 4234 -1041
rect 4238 -1043 4258 -1041
rect 4198 -1045 4258 -1043
rect 4262 -1045 4287 -1041
rect 4198 -1051 4202 -1045
rect 4222 -1051 4226 -1045
rect 4255 -1051 4258 -1045
rect 4211 -1062 4215 -1055
rect 4170 -1066 4204 -1063
rect 4211 -1065 4226 -1062
rect 4222 -1068 4226 -1065
rect 3883 -1079 3887 -1072
rect 4205 -1071 4215 -1070
rect 3790 -1083 3876 -1080
rect 3883 -1082 3898 -1079
rect 3894 -1085 3898 -1082
rect 3877 -1088 3887 -1087
rect 3822 -1091 3887 -1088
rect 3894 -1088 3899 -1085
rect 3943 -1087 3946 -1073
rect 4172 -1074 4215 -1071
rect 4222 -1071 4227 -1068
rect 4271 -1069 4274 -1056
rect 3012 -1095 3058 -1092
rect 3068 -1095 3072 -1092
rect 3040 -1096 3072 -1095
rect 3040 -1098 3048 -1096
rect 3052 -1098 3072 -1096
rect 3021 -1169 3337 -1165
rect 3020 -1184 3164 -1180
rect 3009 -1217 3022 -1213
rect 3026 -1215 3030 -1213
rect 3034 -1215 3050 -1213
rect 3026 -1217 3050 -1215
rect 3019 -1223 3022 -1217
rect 3035 -1243 3038 -1228
rect 3025 -1247 3026 -1243
rect 3035 -1246 3062 -1243
rect 3035 -1262 3038 -1246
rect 3019 -1274 3023 -1267
rect 3009 -1279 3051 -1274
rect 3009 -1280 3025 -1279
rect 3029 -1280 3051 -1279
rect 3059 -1348 3062 -1246
rect 3095 -1286 3098 -1191
rect 3160 -1242 3164 -1184
rect 3186 -1216 3199 -1212
rect 3203 -1214 3207 -1212
rect 3211 -1214 3227 -1212
rect 3203 -1216 3227 -1214
rect 3196 -1222 3199 -1216
rect 3212 -1242 3215 -1227
rect 3160 -1246 3203 -1242
rect 3212 -1245 3255 -1242
rect 3212 -1261 3215 -1245
rect 3196 -1273 3200 -1266
rect 3186 -1278 3228 -1273
rect 3186 -1279 3203 -1278
rect 3207 -1279 3228 -1278
rect 3081 -1327 3086 -1326
rect 3071 -1329 3107 -1327
rect 3111 -1329 3131 -1327
rect 3071 -1331 3131 -1329
rect 3135 -1331 3160 -1327
rect 3071 -1337 3075 -1331
rect 3095 -1337 3099 -1331
rect 3128 -1337 3131 -1331
rect 3084 -1348 3088 -1341
rect 3059 -1352 3077 -1348
rect 3084 -1351 3099 -1348
rect 3095 -1354 3099 -1351
rect 3070 -1360 3088 -1356
rect 3095 -1357 3100 -1354
rect 3144 -1357 3147 -1342
rect 3252 -1352 3255 -1245
rect 3333 -1243 3337 -1169
rect 3361 -1217 3374 -1213
rect 3378 -1215 3382 -1213
rect 3386 -1215 3402 -1213
rect 3378 -1217 3402 -1215
rect 3371 -1223 3374 -1217
rect 3387 -1243 3390 -1228
rect 3333 -1247 3378 -1243
rect 3387 -1246 3436 -1243
rect 3387 -1262 3390 -1246
rect 3371 -1274 3375 -1267
rect 3361 -1279 3403 -1274
rect 3361 -1280 3378 -1279
rect 3382 -1280 3403 -1279
rect 3274 -1331 3279 -1330
rect 3264 -1333 3299 -1331
rect 3303 -1333 3324 -1331
rect 3264 -1335 3324 -1333
rect 3328 -1335 3353 -1331
rect 3264 -1341 3268 -1335
rect 3288 -1341 3292 -1335
rect 3321 -1341 3324 -1335
rect 3277 -1352 3281 -1345
rect 3252 -1356 3270 -1352
rect 3277 -1355 3292 -1352
rect 2924 -1366 2964 -1362
rect 2973 -1365 2998 -1362
rect 3095 -1361 3135 -1357
rect 3144 -1360 3179 -1357
rect 3288 -1358 3292 -1355
rect 2924 -1373 2928 -1366
rect 2901 -1386 2905 -1377
rect 2973 -1381 2976 -1365
rect 3095 -1368 3099 -1361
rect 3072 -1381 3076 -1372
rect 3144 -1376 3147 -1360
rect 3072 -1384 3118 -1381
rect 3128 -1384 3132 -1381
rect 3100 -1386 3132 -1384
rect 2875 -1389 2947 -1386
rect 2957 -1389 2961 -1386
rect 3100 -1387 3110 -1386
rect 2929 -1391 2961 -1389
rect 3114 -1387 3132 -1386
rect 2929 -1392 2939 -1391
rect 2943 -1392 2961 -1391
rect 3176 -1450 3179 -1360
rect 3264 -1364 3281 -1360
rect 3288 -1361 3293 -1358
rect 3337 -1360 3340 -1346
rect 3433 -1348 3436 -1246
rect 3455 -1327 3460 -1326
rect 3445 -1329 3482 -1327
rect 3486 -1329 3505 -1327
rect 3445 -1331 3505 -1329
rect 3509 -1331 3534 -1327
rect 3445 -1337 3449 -1331
rect 3469 -1337 3473 -1331
rect 3502 -1337 3505 -1331
rect 3458 -1348 3462 -1341
rect 3433 -1352 3451 -1348
rect 3458 -1351 3473 -1348
rect 3469 -1354 3473 -1351
rect 3445 -1360 3462 -1356
rect 3469 -1357 3474 -1354
rect 3518 -1356 3521 -1342
rect 3288 -1365 3328 -1361
rect 3337 -1363 3365 -1360
rect 3288 -1372 3292 -1365
rect 3265 -1385 3269 -1376
rect 3337 -1380 3340 -1363
rect 3265 -1388 3311 -1385
rect 3321 -1388 3325 -1385
rect 3293 -1390 3325 -1388
rect 3293 -1391 3303 -1390
rect 3307 -1391 3325 -1390
rect 3362 -1405 3365 -1363
rect 3469 -1361 3509 -1357
rect 3518 -1360 3523 -1356
rect 3469 -1368 3473 -1361
rect 3446 -1381 3450 -1372
rect 3518 -1376 3521 -1360
rect 3446 -1384 3492 -1381
rect 3502 -1384 3506 -1381
rect 3474 -1386 3506 -1384
rect 3474 -1387 3484 -1386
rect 3488 -1387 3506 -1386
rect 3822 -1405 3825 -1091
rect 3894 -1092 3934 -1088
rect 3943 -1091 3948 -1087
rect 3894 -1099 3898 -1092
rect 3871 -1112 3875 -1103
rect 3943 -1107 3946 -1091
rect 3871 -1115 3917 -1112
rect 3927 -1115 3931 -1112
rect 3899 -1116 3931 -1115
rect 3899 -1118 3907 -1116
rect 3911 -1118 3931 -1116
rect 3362 -1408 3825 -1405
rect 4172 -1450 4175 -1074
rect 4222 -1075 4262 -1071
rect 4271 -1075 4277 -1069
rect 4222 -1082 4226 -1075
rect 4199 -1095 4203 -1086
rect 4271 -1090 4274 -1075
rect 4199 -1097 4245 -1095
rect 4255 -1097 4259 -1095
rect 4199 -1098 4259 -1097
rect 4227 -1099 4259 -1098
rect 4227 -1101 4242 -1099
rect 4246 -1101 4259 -1099
rect 3176 -1453 4175 -1450
rect 3667 -1528 3672 -1527
rect 3657 -1530 3705 -1528
rect 3710 -1529 3750 -1528
rect 3710 -1530 3763 -1529
rect 3657 -1532 3763 -1530
rect 3657 -1538 3661 -1532
rect 3681 -1538 3685 -1532
rect 3735 -1533 3763 -1532
rect 3735 -1539 3739 -1533
rect 3759 -1539 3763 -1533
rect 3670 -1549 3674 -1542
rect 3653 -1553 3663 -1549
rect 3670 -1552 3685 -1549
rect 3748 -1550 3752 -1543
rect 3656 -1557 3659 -1553
rect 3681 -1555 3685 -1552
rect 3733 -1554 3741 -1550
rect 3748 -1553 3763 -1550
rect 3656 -1561 3674 -1557
rect 3681 -1558 3686 -1555
rect 3733 -1558 3737 -1554
rect 3759 -1556 3763 -1553
rect 3759 -1558 3764 -1556
rect 3681 -1562 3693 -1558
rect 3733 -1562 3752 -1558
rect 3759 -1561 3771 -1558
rect 3681 -1569 3685 -1562
rect 3658 -1582 3662 -1573
rect 3658 -1585 3687 -1582
rect 3667 -1586 3675 -1585
rect 3667 -1587 3671 -1586
rect 3690 -1652 3693 -1562
rect 3759 -1570 3763 -1561
rect 3736 -1583 3740 -1574
rect 3736 -1585 3765 -1583
rect 3736 -1586 3757 -1585
rect 3747 -1588 3753 -1586
rect 3761 -1586 3765 -1585
rect 3768 -1612 3771 -1561
rect 3696 -1615 3771 -1612
rect 3696 -1644 3700 -1615
rect 3714 -1625 3726 -1623
rect 3731 -1625 3742 -1623
rect 3714 -1627 3742 -1625
rect 3714 -1633 3718 -1627
rect 3738 -1633 3742 -1627
rect 4548 -1629 4561 -1625
rect 4565 -1627 4570 -1625
rect 4574 -1627 4589 -1625
rect 4565 -1629 4589 -1627
rect 4558 -1635 4561 -1629
rect 3727 -1644 3731 -1637
rect 4012 -1638 4017 -1637
rect 4002 -1640 4051 -1638
rect 4055 -1639 4095 -1638
rect 4055 -1640 4108 -1639
rect 4002 -1642 4108 -1640
rect 3696 -1648 3720 -1644
rect 3727 -1647 3742 -1644
rect 3738 -1650 3742 -1647
rect 4002 -1648 4006 -1642
rect 4026 -1648 4030 -1642
rect 3690 -1656 3731 -1652
rect 3738 -1654 3744 -1650
rect 4080 -1643 4108 -1642
rect 4080 -1649 4084 -1643
rect 4104 -1649 4108 -1643
rect 3738 -1664 3742 -1654
rect 4015 -1659 4019 -1652
rect 3982 -1663 4008 -1659
rect 4015 -1662 4030 -1659
rect 4093 -1660 4097 -1653
rect 4574 -1655 4577 -1640
rect 4897 -1655 4901 -1027
rect 5032 -1028 5072 -1024
rect 5081 -1027 5242 -1024
rect 5032 -1035 5036 -1028
rect 5009 -1048 5013 -1039
rect 5081 -1043 5084 -1027
rect 5232 -1028 5242 -1027
rect 5249 -1025 5254 -1022
rect 5298 -1025 5301 -1010
rect 5249 -1029 5289 -1025
rect 5298 -1028 5329 -1025
rect 5249 -1036 5253 -1029
rect 5009 -1051 5055 -1048
rect 5065 -1051 5069 -1048
rect 5037 -1053 5069 -1051
rect 5226 -1049 5230 -1040
rect 5298 -1044 5301 -1028
rect 5226 -1052 5272 -1049
rect 5282 -1052 5286 -1049
rect 5037 -1054 5046 -1053
rect 5050 -1054 5069 -1053
rect 5254 -1054 5286 -1052
rect 5254 -1055 5258 -1054
rect 5262 -1055 5286 -1054
rect 4490 -1659 4565 -1655
rect 4574 -1659 4901 -1655
rect 3715 -1677 3719 -1668
rect 3715 -1680 3744 -1677
rect 3726 -1681 3734 -1680
rect 3726 -1682 3729 -1681
rect 3733 -1682 3734 -1681
rect 3677 -1772 3682 -1771
rect 3667 -1774 3710 -1772
rect 3714 -1773 3760 -1772
rect 3714 -1774 3773 -1773
rect 3667 -1776 3773 -1774
rect 3667 -1782 3671 -1776
rect 3691 -1782 3695 -1776
rect 3745 -1777 3773 -1776
rect 3745 -1783 3749 -1777
rect 3769 -1783 3773 -1777
rect 3680 -1793 3684 -1786
rect 3663 -1797 3673 -1793
rect 3680 -1796 3695 -1793
rect 3758 -1794 3762 -1787
rect 3666 -1801 3669 -1797
rect 3691 -1799 3695 -1796
rect 3743 -1798 3751 -1794
rect 3758 -1797 3773 -1794
rect 3666 -1805 3684 -1801
rect 3691 -1802 3696 -1799
rect 3743 -1802 3747 -1798
rect 3769 -1800 3773 -1797
rect 3769 -1802 3774 -1800
rect 3691 -1806 3703 -1802
rect 3743 -1806 3762 -1802
rect 3769 -1805 3781 -1802
rect 3691 -1813 3695 -1806
rect 3668 -1826 3672 -1817
rect 3668 -1829 3697 -1826
rect 3677 -1830 3684 -1829
rect 3677 -1831 3678 -1830
rect 3682 -1831 3684 -1830
rect 3700 -1896 3703 -1806
rect 3769 -1814 3773 -1805
rect 3746 -1827 3750 -1818
rect 3746 -1830 3775 -1827
rect 3757 -1831 3763 -1830
rect 3757 -1832 3759 -1831
rect 3778 -1856 3781 -1805
rect 3706 -1859 3781 -1856
rect 3706 -1888 3710 -1859
rect 3738 -1866 3741 -1864
rect 3734 -1867 3741 -1866
rect 3724 -1871 3752 -1867
rect 3724 -1877 3728 -1871
rect 3748 -1877 3752 -1871
rect 3737 -1888 3741 -1881
rect 3706 -1892 3730 -1888
rect 3737 -1891 3752 -1888
rect 3748 -1894 3752 -1891
rect 3982 -1894 3986 -1663
rect 4001 -1667 4004 -1663
rect 4026 -1665 4030 -1662
rect 4078 -1664 4086 -1660
rect 4093 -1663 4108 -1660
rect 4001 -1671 4019 -1667
rect 4026 -1668 4031 -1665
rect 4078 -1668 4082 -1664
rect 4104 -1666 4108 -1663
rect 4104 -1668 4109 -1666
rect 4026 -1672 4038 -1668
rect 4078 -1672 4097 -1668
rect 4104 -1671 4116 -1668
rect 4026 -1679 4030 -1672
rect 4003 -1692 4007 -1683
rect 4003 -1695 4032 -1692
rect 4012 -1696 4019 -1695
rect 4012 -1697 4015 -1696
rect 4035 -1762 4038 -1672
rect 4104 -1680 4108 -1671
rect 4081 -1693 4085 -1684
rect 4081 -1696 4110 -1693
rect 4092 -1697 4098 -1696
rect 4092 -1698 4094 -1697
rect 4113 -1722 4116 -1671
rect 4041 -1725 4116 -1722
rect 4041 -1754 4045 -1725
rect 4069 -1733 4073 -1732
rect 4059 -1737 4087 -1733
rect 4059 -1743 4063 -1737
rect 4083 -1743 4087 -1737
rect 4072 -1754 4076 -1747
rect 4041 -1758 4065 -1754
rect 4072 -1757 4087 -1754
rect 4083 -1760 4087 -1757
rect 4490 -1760 4494 -1659
rect 4574 -1674 4577 -1659
rect 4558 -1686 4562 -1679
rect 4548 -1691 4590 -1686
rect 4548 -1692 4565 -1691
rect 4569 -1692 4590 -1691
rect 4035 -1766 4076 -1762
rect 4083 -1764 4494 -1760
rect 4083 -1774 4087 -1764
rect 4060 -1787 4064 -1778
rect 4060 -1790 4089 -1787
rect 4071 -1791 4079 -1790
rect 4071 -1792 4073 -1791
rect 4077 -1792 4079 -1791
rect 3700 -1900 3741 -1896
rect 3748 -1898 3986 -1894
rect 3748 -1908 3752 -1898
rect 3725 -1921 3729 -1912
rect 3725 -1924 3754 -1921
rect 3736 -1925 3744 -1924
rect 3736 -1926 3738 -1925
rect 3742 -1926 3744 -1925
<< metal2 >>
rect 3024 837 5243 841
rect 3024 835 5239 837
rect 3024 732 3030 835
rect 3151 755 3360 759
rect 2695 728 3045 732
rect 2695 466 2699 728
rect 1196 462 2699 466
rect 2826 685 3000 689
rect 964 250 1072 254
rect 964 231 968 250
rect 1068 235 1072 250
rect 1068 231 1077 235
rect 937 227 968 231
rect 937 46 941 227
rect 964 215 968 227
rect 1196 226 1200 462
rect 1307 427 1311 462
rect 1307 423 1328 427
rect 2826 422 2830 685
rect 2996 667 3000 685
rect 3042 630 3045 728
rect 3042 626 3043 630
rect 2973 519 3096 523
rect 2973 501 2977 519
rect 3092 512 3096 519
rect 2889 497 2977 501
rect 2915 422 2918 457
rect 2826 419 2918 422
rect 1281 387 1348 389
rect 1281 386 1352 387
rect 2826 373 2830 419
rect 2974 381 2977 497
rect 3120 457 3122 461
rect 3120 421 3124 457
rect 3151 421 3155 755
rect 3120 417 3155 421
rect 3163 470 3288 473
rect 2974 377 3004 381
rect 2826 369 2849 373
rect 2993 369 3004 373
rect 3163 372 3166 470
rect 3285 435 3288 470
rect 3285 431 3300 435
rect 3243 396 3244 398
rect 3239 395 3244 396
rect 3318 395 3322 396
rect 3239 391 3322 395
rect 3092 369 3166 372
rect 1165 222 1200 226
rect 1411 356 1417 360
rect 1411 158 1415 356
rect 1524 160 1528 362
rect 1633 358 1644 362
rect 1757 359 1764 363
rect 1633 160 1637 358
rect 1757 161 1762 359
rect 1941 162 1946 364
rect 2030 359 2035 363
rect 2054 362 2057 366
rect 2141 362 2151 366
rect 2166 362 2173 366
rect 2031 223 2035 359
rect 2147 250 2151 362
rect 2256 360 2264 364
rect 2288 363 2296 367
rect 2260 275 2264 360
rect 2993 285 2997 369
rect 3352 285 3356 755
rect 2993 281 3356 285
rect 3514 735 3757 739
rect 3514 275 3518 735
rect 3566 701 3740 705
rect 3566 438 3570 701
rect 3736 683 3740 701
rect 3753 693 3757 735
rect 3782 646 3785 835
rect 4561 834 4565 835
rect 3891 771 4100 775
rect 3782 642 3783 646
rect 3713 535 3836 539
rect 3713 517 3717 535
rect 3832 528 3836 535
rect 3629 513 3717 517
rect 3655 438 3658 473
rect 3566 435 3658 438
rect 3550 393 3552 397
rect 2260 271 3519 275
rect 3550 255 3554 393
rect 3566 389 3570 435
rect 3714 397 3717 513
rect 3860 473 3862 477
rect 3860 437 3864 473
rect 3891 437 3895 771
rect 3860 433 3895 437
rect 3903 486 4028 489
rect 3714 393 3744 397
rect 3566 385 3589 389
rect 3733 385 3744 389
rect 3903 388 3906 486
rect 4025 451 4028 486
rect 4025 447 4040 451
rect 3990 412 4045 416
rect 3832 385 3906 388
rect 3733 301 3737 385
rect 4092 301 4096 771
rect 3733 297 4096 301
rect 4312 745 4538 749
rect 2147 246 3201 250
rect 3197 231 3201 246
rect 4312 231 4316 745
rect 4345 712 4519 716
rect 4345 449 4349 712
rect 4515 694 4519 712
rect 4534 703 4538 745
rect 4561 657 4564 834
rect 4670 782 5585 786
rect 4561 653 4562 657
rect 4492 546 4615 550
rect 4492 528 4496 546
rect 4611 539 4615 546
rect 4408 524 4496 528
rect 4434 449 4437 484
rect 4345 446 4437 449
rect 4327 404 4330 408
rect 4327 243 4332 404
rect 4345 400 4349 446
rect 4493 408 4496 524
rect 4639 484 4641 488
rect 4639 448 4643 484
rect 4670 448 4674 782
rect 4639 444 4674 448
rect 4682 497 4807 500
rect 4493 404 4523 408
rect 4345 396 4368 400
rect 4512 396 4523 400
rect 4682 399 4685 497
rect 4804 462 4807 497
rect 4804 458 4819 462
rect 4758 419 4762 423
rect 4837 419 4841 422
rect 4758 416 4841 419
rect 4611 396 4685 399
rect 4512 312 4516 396
rect 4920 312 4924 782
rect 4512 308 4924 312
rect 5000 726 5215 730
rect 4327 240 4328 243
rect 3197 227 4316 231
rect 5000 223 5004 726
rect 5025 706 5199 710
rect 5025 443 5029 706
rect 5195 688 5199 706
rect 5211 697 5215 726
rect 5241 688 5244 690
rect 5241 685 5323 688
rect 5241 651 5244 685
rect 5241 647 5242 651
rect 5172 540 5295 544
rect 5172 522 5176 540
rect 5291 533 5295 540
rect 5088 518 5176 522
rect 5114 443 5117 478
rect 5025 440 5117 443
rect 5025 394 5029 440
rect 5173 402 5176 518
rect 5320 489 5323 685
rect 5362 491 5487 494
rect 5320 485 5321 489
rect 5173 398 5203 402
rect 5025 390 5048 394
rect 5362 393 5365 491
rect 5484 456 5487 491
rect 5484 452 5499 456
rect 5442 413 5446 417
rect 5517 413 5521 416
rect 5442 410 5521 413
rect 5291 390 5365 393
rect 5581 356 5585 782
rect 5525 352 5585 356
rect 2031 219 5004 223
rect 1411 154 1420 158
rect 1524 156 1531 160
rect 1633 156 1647 160
rect 1757 157 1767 161
rect 1941 158 1949 162
rect 1049 131 1076 135
rect 937 42 1078 46
rect 1411 -19 1415 154
rect 1524 60 1528 156
rect 1524 56 1553 60
rect 1549 -17 1553 56
rect 1633 53 1637 156
rect 1757 64 1762 157
rect 1757 59 1788 64
rect 1633 49 1668 53
rect 1664 -17 1668 49
rect 1783 -16 1788 59
rect 1941 -15 1946 158
rect 2037 157 2043 161
rect 2054 160 2060 164
rect 2147 158 2157 163
rect 2166 160 2176 164
rect 2265 159 2278 163
rect 2288 161 2296 165
rect 2384 160 2393 164
rect 2039 71 2043 157
rect 2152 82 2157 158
rect 2274 91 2278 159
rect 2389 101 2393 160
rect 2389 97 2540 101
rect 2274 87 2529 91
rect 2152 77 2519 82
rect 2039 67 2505 71
rect 1411 -23 1445 -19
rect 1549 -21 1556 -17
rect 1664 -21 1672 -17
rect 1783 -20 1792 -16
rect 1941 -19 1974 -15
rect 2078 -17 2085 -13
rect 2198 -17 2201 -13
rect 2320 -16 2323 -12
rect 2062 -72 2066 -65
rect 2182 -66 2186 -54
rect 2182 -70 2456 -66
rect 1688 -76 2066 -72
rect 1688 -160 1692 -76
rect 1688 -164 1712 -160
rect 1816 -165 1819 -161
rect 1956 -165 1963 -161
rect 1816 -241 1820 -165
rect 1956 -225 1959 -165
rect 2287 -225 2290 -208
rect 1956 -228 2290 -225
rect 2452 -241 2456 -70
rect 1816 -245 2456 -241
rect 2501 -731 2505 67
rect 2514 -534 2519 77
rect 2514 -692 2518 -534
rect 2525 -678 2529 87
rect 2536 -665 2540 97
rect 2743 1 3575 5
rect 2536 -669 2707 -665
rect 2525 -682 2708 -678
rect 2514 -696 2710 -692
rect 2501 -735 2713 -731
rect 2743 -933 2747 1
rect 3646 -1 3654 4
rect 3646 -49 3650 -1
rect 3646 -53 4422 -49
rect 3750 -91 3858 -86
rect 3750 -96 3755 -91
rect 3676 -100 3755 -96
rect 3675 -101 3755 -100
rect 3853 -123 3858 -91
rect 3853 -128 3872 -123
rect 3533 -275 3588 -271
rect 2769 -534 3306 -530
rect 2768 -555 3145 -551
rect 2768 -571 2958 -567
rect 2769 -613 2830 -611
rect 2769 -616 2775 -613
rect 2779 -616 2830 -613
rect 2956 -612 2960 -571
rect 3143 -611 3147 -555
rect 2956 -614 2996 -612
rect 2956 -616 2974 -614
rect 2971 -617 2974 -616
rect 2978 -616 2996 -614
rect 3143 -613 3171 -611
rect 3143 -615 3154 -613
rect 3151 -616 3154 -615
rect 2978 -617 2983 -616
rect 3158 -615 3171 -613
rect 3304 -612 3308 -534
rect 3304 -614 3348 -612
rect 3158 -616 3163 -615
rect 3304 -616 3332 -614
rect 3330 -617 3332 -616
rect 3336 -616 3348 -614
rect 3336 -617 3339 -616
rect 2834 -654 2838 -652
rect 3001 -654 3006 -652
rect 3178 -654 3183 -651
rect 3353 -654 3357 -652
rect 2834 -658 3357 -654
rect 2810 -669 3389 -665
rect 2796 -682 3186 -678
rect 2777 -696 3011 -692
rect 3007 -725 3011 -696
rect 3007 -727 3041 -725
rect 3007 -729 3021 -727
rect 2816 -731 2870 -730
rect 2762 -732 2870 -731
rect 2762 -734 2842 -732
rect 2762 -735 2816 -734
rect 2846 -734 2870 -732
rect 3025 -729 3041 -727
rect 3127 -729 3146 -725
rect 2960 -821 2984 -817
rect 3089 -873 3103 -869
rect 3099 -933 3103 -873
rect 2743 -937 3103 -933
rect 3142 -961 3146 -729
rect 3182 -729 3186 -682
rect 3385 -725 3389 -669
rect 3533 -725 3537 -275
rect 3659 -277 3667 -272
rect 3659 -325 3663 -277
rect 3659 -329 3955 -325
rect 3860 -530 3866 -529
rect 3860 -538 3866 -537
rect 3723 -615 3842 -612
rect 3723 -657 3727 -615
rect 3838 -630 3842 -615
rect 3862 -622 3866 -538
rect 3723 -661 3746 -657
rect 3885 -672 3886 -668
rect 3751 -701 3756 -697
rect 3875 -701 3879 -693
rect 3751 -704 3879 -701
rect 3885 -708 3888 -672
rect 3385 -729 3415 -725
rect 3501 -729 3537 -725
rect 3566 -712 3888 -708
rect 3182 -731 3234 -729
rect 3182 -733 3210 -731
rect 3214 -733 3234 -731
rect 3329 -734 3346 -730
rect 3342 -894 3346 -734
rect 3385 -761 3389 -729
rect 3566 -761 3570 -712
rect 3385 -765 3570 -761
rect 3342 -898 3849 -894
rect 3951 -901 3955 -329
rect 4103 -550 4109 -549
rect 4103 -558 4109 -557
rect 3971 -616 4090 -613
rect 3971 -658 3975 -616
rect 4086 -631 4090 -616
rect 4105 -623 4109 -558
rect 4345 -567 4351 -566
rect 4345 -575 4351 -574
rect 3971 -662 3994 -658
rect 4015 -662 4056 -658
rect 4053 -779 4056 -662
rect 4132 -668 4136 -582
rect 4214 -607 4333 -604
rect 4214 -649 4218 -607
rect 4329 -622 4333 -607
rect 4346 -614 4350 -575
rect 4214 -653 4237 -649
rect 4375 -659 4379 -593
rect 4375 -663 4377 -659
rect 4132 -672 4134 -668
rect 4244 -694 4248 -689
rect 4369 -694 4373 -685
rect 4244 -698 4373 -694
rect 4053 -783 4070 -779
rect 3938 -905 3955 -901
rect 4224 -803 4290 -799
rect 4224 -961 4228 -803
rect 4418 -806 4422 -53
rect 4483 -602 4602 -599
rect 4483 -644 4487 -602
rect 4598 -617 4602 -602
rect 4618 -609 4622 -566
rect 4483 -648 4506 -644
rect 4645 -654 4648 -595
rect 4645 -658 4646 -654
rect 4380 -810 4422 -806
rect 3142 -965 4228 -961
rect 3093 -1071 3128 -1067
rect 3124 -1153 3128 -1071
rect 4285 -1075 4309 -1069
rect 3952 -1091 3973 -1087
rect 2773 -1157 3128 -1153
rect 2773 -1690 2777 -1157
rect 2983 -1169 3015 -1165
rect 2983 -1184 3013 -1180
rect 2986 -1247 3021 -1243
rect 2858 -1288 2862 -1282
rect 3025 -1288 3029 -1283
rect 2858 -1290 3094 -1288
rect 3203 -1288 3207 -1282
rect 3378 -1288 3382 -1283
rect 3098 -1290 3382 -1288
rect 2858 -1292 3382 -1290
rect 3054 -1358 3066 -1356
rect 2884 -1365 2896 -1361
rect 3041 -1360 3066 -1358
rect 3070 -1360 3071 -1356
rect 3041 -1364 3057 -1360
rect 3251 -1364 3260 -1360
rect 3410 -1356 3416 -1355
rect 3410 -1360 3439 -1356
rect 3527 -1360 3623 -1356
rect 3410 -1361 3442 -1360
rect 2884 -1376 2888 -1365
rect 3232 -1370 3254 -1364
rect 2872 -1382 2888 -1376
rect 3619 -1549 3623 -1360
rect 3619 -1553 3647 -1549
rect 3718 -1555 3726 -1550
rect 3718 -1602 3722 -1555
rect 3969 -1602 3973 -1091
rect 3718 -1606 3973 -1602
rect 3768 -1607 3771 -1606
rect 3977 -1630 4069 -1625
rect 3977 -1650 3982 -1630
rect 3748 -1654 3982 -1650
rect 3747 -1655 3982 -1654
rect 4064 -1660 4069 -1630
rect 4064 -1665 4071 -1660
rect 2773 -1694 3633 -1690
rect 3629 -1793 3633 -1694
rect 3629 -1797 3657 -1793
rect 3728 -1799 3736 -1794
rect 3728 -1846 3732 -1799
rect 4303 -1846 4309 -1075
rect 3728 -1850 4309 -1846
rect 3778 -1851 3781 -1850
<< metal3 >>
rect 2282 367 2289 368
rect 2049 366 2055 367
rect 2049 362 2050 366
rect 2054 362 2055 366
rect 2049 164 2055 362
rect 2049 160 2050 164
rect 2054 160 2055 164
rect 2049 91 2055 160
rect 2160 366 2167 367
rect 2160 362 2161 366
rect 2166 362 2167 366
rect 2160 164 2167 362
rect 2160 160 2161 164
rect 2166 160 2167 164
rect 2160 98 2167 160
rect 2282 363 2283 367
rect 2288 363 2289 367
rect 2282 165 2289 363
rect 2282 161 2283 165
rect 2288 161 2289 165
rect 2282 102 2289 161
rect 2160 91 2199 98
rect 2282 95 2321 102
rect 2049 85 2079 91
rect 2073 -13 2079 85
rect 2073 -17 2074 -13
rect 2078 -17 2079 -13
rect 2073 -18 2079 -17
rect 2192 -13 2199 91
rect 2192 -17 2194 -13
rect 2198 -17 2199 -13
rect 2314 -12 2321 95
rect 2314 -16 2315 -12
rect 2320 -16 2321 -12
rect 2314 -17 2321 -16
rect 2192 -18 2199 -17
rect 3304 -530 3867 -529
rect 3304 -534 3306 -530
rect 3310 -534 3860 -530
rect 3304 -535 3860 -534
rect 3859 -537 3860 -535
rect 3866 -537 3867 -530
rect 3859 -538 3867 -537
rect 4101 -550 4110 -549
rect 3143 -551 4103 -550
rect 3143 -555 3145 -551
rect 3149 -555 4103 -551
rect 3143 -556 4103 -555
rect 4102 -557 4103 -556
rect 4109 -557 4110 -550
rect 4102 -558 4110 -557
rect 4616 -561 4624 -560
rect 4616 -566 4618 -561
rect 4623 -566 4689 -561
rect 2956 -567 4352 -566
rect 4616 -567 4689 -566
rect 2956 -571 2958 -567
rect 2962 -571 4345 -567
rect 2956 -572 4345 -571
rect 4343 -573 4345 -572
rect 4344 -574 4345 -573
rect 4351 -574 4352 -567
rect 4344 -575 4352 -574
rect 2773 -613 2781 -611
rect 2773 -618 2775 -613
rect 2779 -618 2781 -613
rect 2972 -614 2980 -612
rect 2774 -1376 2780 -618
rect 2972 -619 2974 -614
rect 2978 -619 2980 -614
rect 3152 -613 3160 -611
rect 3152 -618 3154 -613
rect 3158 -618 3160 -613
rect 3330 -614 3338 -612
rect 2973 -1301 2979 -619
rect 2973 -1307 3034 -1301
rect 3028 -1353 3034 -1307
rect 3153 -1305 3159 -618
rect 3330 -619 3332 -614
rect 3336 -619 3338 -614
rect 3331 -1298 3337 -619
rect 3331 -1304 3407 -1298
rect 3153 -1311 3230 -1305
rect 3028 -1357 3035 -1353
rect 3028 -1358 3043 -1357
rect 3028 -1364 3036 -1358
rect 3041 -1364 3043 -1358
rect 3035 -1366 3043 -1364
rect 3224 -1360 3230 -1311
rect 3401 -1351 3407 -1304
rect 3401 -1355 3416 -1351
rect 3224 -1364 3234 -1360
rect 3401 -1361 3405 -1355
rect 3410 -1361 3416 -1355
rect 3401 -1363 3416 -1361
rect 3224 -1370 3227 -1364
rect 3232 -1370 3234 -1364
rect 3226 -1372 3234 -1370
rect 2866 -1376 2874 -1375
rect 2774 -1382 2867 -1376
rect 2872 -1382 2874 -1376
rect 2840 -1428 2846 -1382
rect 2866 -1384 2874 -1382
rect 4683 -1428 4689 -567
rect 2840 -1434 4689 -1428
<< ntransistor >>
rect 2988 611 2990 616
rect 3007 611 3009 616
rect 3032 611 3034 616
rect 3051 611 3053 616
rect 3728 627 3730 632
rect 3747 627 3749 632
rect 3772 627 3774 632
rect 3791 627 3793 632
rect 4507 638 4509 643
rect 4526 638 4528 643
rect 4551 638 4553 643
rect 4570 638 4572 643
rect 1265 399 1268 408
rect 1276 399 1279 408
rect 1088 289 1091 298
rect 1099 289 1102 298
rect 1146 285 1149 290
rect 2862 445 2864 450
rect 2881 445 2883 450
rect 2906 445 2908 450
rect 2925 445 2927 450
rect 3067 449 3069 454
rect 3086 449 3088 454
rect 3111 449 3113 454
rect 3130 449 3132 454
rect 1343 398 1346 407
rect 1354 398 1357 407
rect 1322 304 1325 313
rect 1333 304 1336 313
rect 1090 206 1093 215
rect 1101 206 1104 215
rect 1148 202 1151 207
rect 989 191 992 196
rect 990 94 993 99
rect 1088 106 1091 115
rect 1099 106 1102 115
rect 1146 102 1149 107
rect 1089 17 1092 26
rect 1100 17 1103 26
rect 1147 13 1150 18
rect 1429 339 1432 348
rect 1440 339 1443 348
rect 1540 341 1543 350
rect 1551 341 1554 350
rect 1487 335 1490 340
rect 1598 337 1601 342
rect 1656 341 1659 350
rect 1667 341 1670 350
rect 1776 342 1779 351
rect 1787 342 1790 351
rect 1958 343 1961 352
rect 1969 343 1972 352
rect 2069 345 2072 354
rect 2080 345 2083 354
rect 1714 337 1717 342
rect 1834 338 1837 343
rect 2016 339 2019 344
rect 2127 341 2130 346
rect 2185 345 2188 354
rect 2196 345 2199 354
rect 2305 346 2308 355
rect 2316 346 2319 355
rect 2862 352 2865 361
rect 2873 352 2876 361
rect 2920 348 2923 353
rect 3017 352 3020 361
rect 3028 352 3031 361
rect 3075 348 3078 353
rect 2243 341 2246 346
rect 2363 342 2366 347
rect 3235 407 3238 416
rect 3246 407 3249 416
rect 3602 461 3604 466
rect 3621 461 3623 466
rect 3646 461 3648 466
rect 3665 461 3667 466
rect 3807 465 3809 470
rect 3826 465 3828 470
rect 3851 465 3853 470
rect 3870 465 3872 470
rect 5187 632 5189 637
rect 5206 632 5208 637
rect 5231 632 5233 637
rect 5250 632 5252 637
rect 3313 406 3316 415
rect 3324 406 3327 415
rect 3602 368 3605 377
rect 3613 368 3616 377
rect 3660 364 3663 369
rect 3757 368 3760 377
rect 3768 368 3771 377
rect 3815 364 3818 369
rect 3975 423 3978 432
rect 3986 423 3989 432
rect 4381 472 4383 477
rect 4400 472 4402 477
rect 4425 472 4427 477
rect 4444 472 4446 477
rect 4586 476 4588 481
rect 4605 476 4607 481
rect 4630 476 4632 481
rect 4649 476 4651 481
rect 4053 422 4056 431
rect 4064 422 4067 431
rect 4381 379 4384 388
rect 4392 379 4395 388
rect 4439 375 4442 380
rect 4536 379 4539 388
rect 4547 379 4550 388
rect 4594 375 4597 380
rect 3292 312 3295 321
rect 3303 312 3306 321
rect 4032 328 4035 337
rect 4043 328 4046 337
rect 4754 434 4757 443
rect 4765 434 4768 443
rect 5061 466 5063 471
rect 5080 466 5082 471
rect 5105 466 5107 471
rect 5124 466 5126 471
rect 4832 433 4835 442
rect 4843 433 4846 442
rect 5266 470 5268 475
rect 5285 470 5287 475
rect 5310 470 5312 475
rect 5329 470 5331 475
rect 5061 373 5064 382
rect 5072 373 5075 382
rect 5119 369 5122 374
rect 5216 373 5219 382
rect 5227 373 5230 382
rect 5274 369 5277 374
rect 5434 428 5437 437
rect 5445 428 5448 437
rect 5512 427 5515 436
rect 5523 427 5526 436
rect 4811 339 4814 348
rect 4822 339 4825 348
rect 5491 333 5494 342
rect 5502 333 5505 342
rect 1432 137 1435 146
rect 1443 137 1446 146
rect 1543 139 1546 148
rect 1554 139 1557 148
rect 1490 133 1493 138
rect 1601 135 1604 140
rect 1659 139 1662 148
rect 1670 139 1673 148
rect 1779 140 1782 149
rect 1790 140 1793 149
rect 1961 141 1964 150
rect 1972 141 1975 150
rect 2072 143 2075 152
rect 2083 143 2086 152
rect 1717 135 1720 140
rect 1837 136 1840 141
rect 2019 137 2022 142
rect 2130 139 2133 144
rect 2188 143 2191 152
rect 2199 143 2202 152
rect 2308 144 2311 153
rect 2319 144 2322 153
rect 2246 139 2249 144
rect 2366 140 2369 145
rect 1457 -40 1460 -31
rect 1468 -40 1471 -31
rect 1568 -38 1571 -29
rect 1579 -38 1582 -29
rect 1515 -44 1518 -39
rect 1626 -42 1629 -37
rect 1684 -38 1687 -29
rect 1695 -38 1698 -29
rect 1804 -37 1807 -28
rect 1815 -37 1818 -28
rect 1986 -36 1989 -27
rect 1997 -36 2000 -27
rect 2097 -34 2100 -25
rect 2108 -34 2111 -25
rect 1742 -42 1745 -37
rect 1862 -41 1865 -36
rect 2044 -40 2047 -35
rect 2155 -38 2158 -33
rect 2213 -34 2216 -25
rect 2224 -34 2227 -25
rect 2333 -33 2336 -24
rect 2344 -33 2347 -24
rect 2271 -38 2274 -33
rect 2391 -37 2394 -32
rect 1724 -181 1727 -172
rect 1735 -181 1738 -172
rect 1782 -185 1785 -180
rect 1842 -182 1845 -173
rect 1853 -182 1856 -173
rect 1900 -186 1903 -181
rect 1975 -182 1978 -173
rect 1986 -182 1989 -173
rect 2033 -186 2036 -181
rect 2094 -183 2097 -174
rect 2105 -183 2108 -174
rect 2152 -187 2155 -182
rect 3592 -24 3595 -15
rect 3603 -24 3606 -15
rect 3670 -25 3673 -16
rect 3681 -25 3684 -16
rect 3649 -119 3652 -110
rect 3660 -119 3663 -110
rect 3810 -151 3813 -142
rect 3821 -151 3824 -142
rect 3605 -300 3608 -291
rect 3616 -300 3619 -291
rect 3888 -152 3891 -143
rect 3899 -152 3902 -143
rect 3867 -246 3870 -237
rect 3878 -246 3881 -237
rect 4104 -192 4107 -187
rect 3683 -301 3686 -292
rect 3694 -301 3697 -292
rect 3662 -395 3665 -386
rect 3673 -395 3676 -386
rect 2837 -636 2840 -631
rect 3002 -636 3005 -631
rect 3179 -635 3182 -630
rect 3354 -636 3357 -631
rect 3752 -681 3755 -676
rect 2882 -751 2885 -742
rect 2893 -751 2896 -742
rect 3053 -746 3056 -737
rect 3064 -746 3067 -737
rect 3111 -750 3114 -745
rect 3246 -750 3249 -741
rect 3257 -750 3260 -741
rect 3427 -746 3430 -737
rect 3438 -746 3441 -737
rect 2940 -755 2943 -750
rect 3304 -754 3307 -749
rect 3485 -750 3488 -745
rect 3014 -890 3017 -881
rect 3025 -890 3028 -881
rect 3072 -894 3075 -889
rect 3018 -1088 3021 -1079
rect 3029 -1088 3032 -1079
rect 3076 -1092 3079 -1087
rect 3831 -686 3833 -681
rect 3850 -686 3852 -681
rect 3875 -686 3877 -681
rect 3894 -686 3896 -681
rect 4000 -682 4003 -677
rect 4079 -687 4081 -682
rect 4098 -687 4100 -682
rect 4123 -687 4125 -682
rect 4142 -687 4144 -682
rect 4243 -673 4246 -668
rect 4322 -678 4324 -673
rect 4341 -678 4343 -673
rect 4366 -678 4368 -673
rect 4385 -678 4387 -673
rect 4512 -668 4515 -663
rect 4591 -673 4593 -668
rect 4610 -673 4612 -668
rect 4635 -673 4637 -668
rect 4654 -673 4656 -668
rect 4085 -807 4088 -798
rect 4096 -807 4099 -798
rect 4143 -811 4146 -806
rect 4305 -827 4308 -818
rect 4316 -827 4319 -818
rect 4461 -819 4464 -810
rect 4472 -819 4475 -810
rect 4519 -823 4522 -818
rect 4363 -831 4366 -826
rect 3864 -922 3867 -913
rect 3875 -922 3878 -913
rect 3922 -926 3925 -921
rect 3877 -1108 3880 -1099
rect 3888 -1108 3891 -1099
rect 3935 -1112 3938 -1107
rect 4205 -1091 4208 -1082
rect 4216 -1091 4219 -1082
rect 4263 -1095 4266 -1090
rect 2862 -1267 2865 -1262
rect 3027 -1267 3030 -1262
rect 3204 -1266 3207 -1261
rect 3379 -1267 3382 -1262
rect 2907 -1382 2910 -1373
rect 2918 -1382 2921 -1373
rect 3078 -1377 3081 -1368
rect 3089 -1377 3092 -1368
rect 3136 -1381 3139 -1376
rect 3271 -1381 3274 -1372
rect 3282 -1381 3285 -1372
rect 3452 -1377 3455 -1368
rect 3463 -1377 3466 -1368
rect 2965 -1386 2968 -1381
rect 3329 -1385 3332 -1380
rect 3510 -1381 3513 -1376
rect 3664 -1578 3667 -1569
rect 3675 -1578 3678 -1569
rect 3742 -1579 3745 -1570
rect 3753 -1579 3756 -1570
rect 5015 -1044 5018 -1035
rect 5026 -1044 5029 -1035
rect 5073 -1048 5076 -1043
rect 5232 -1045 5235 -1036
rect 5243 -1045 5246 -1036
rect 5290 -1049 5293 -1044
rect 3721 -1673 3724 -1664
rect 3732 -1673 3735 -1664
rect 4009 -1688 4012 -1679
rect 4020 -1688 4023 -1679
rect 3674 -1822 3677 -1813
rect 3685 -1822 3688 -1813
rect 4566 -1679 4569 -1674
rect 4087 -1689 4090 -1680
rect 4098 -1689 4101 -1680
rect 4066 -1783 4069 -1774
rect 4077 -1783 4080 -1774
rect 3752 -1823 3755 -1814
rect 3763 -1823 3766 -1814
rect 3731 -1917 3734 -1908
rect 3742 -1917 3745 -1908
<< ptransistor >>
rect 2988 642 2990 647
rect 3007 642 3009 647
rect 3032 642 3034 647
rect 3051 642 3053 647
rect 3728 658 3730 663
rect 3747 658 3749 663
rect 3772 658 3774 663
rect 3791 658 3793 663
rect 4507 669 4509 674
rect 4526 669 4528 674
rect 4551 669 4553 674
rect 4570 669 4572 674
rect 1265 432 1268 439
rect 1276 432 1279 439
rect 1088 322 1091 329
rect 1099 322 1102 329
rect 1146 324 1149 329
rect 1343 431 1346 438
rect 1354 431 1357 438
rect 2862 476 2864 481
rect 2881 476 2883 481
rect 2906 476 2908 481
rect 2925 476 2927 481
rect 3067 480 3069 485
rect 3086 480 3088 485
rect 3111 480 3113 485
rect 3130 480 3132 485
rect 3235 440 3238 447
rect 3246 440 3249 447
rect 1322 337 1325 344
rect 1333 337 1336 344
rect 1090 239 1093 246
rect 1101 239 1104 246
rect 1148 241 1151 246
rect 989 230 992 235
rect 990 133 993 138
rect 1088 139 1091 146
rect 1099 139 1102 146
rect 1146 141 1149 146
rect 1089 50 1092 57
rect 1100 50 1103 57
rect 1147 52 1150 57
rect 1429 372 1432 379
rect 1440 372 1443 379
rect 1487 374 1490 379
rect 1540 374 1543 381
rect 1551 374 1554 381
rect 1598 376 1601 381
rect 1656 374 1659 381
rect 1667 374 1670 381
rect 1714 376 1717 381
rect 1776 375 1779 382
rect 1787 375 1790 382
rect 1834 377 1837 382
rect 1958 376 1961 383
rect 1969 376 1972 383
rect 2016 378 2019 383
rect 2069 378 2072 385
rect 2080 378 2083 385
rect 2127 380 2130 385
rect 2185 378 2188 385
rect 2196 378 2199 385
rect 2243 380 2246 385
rect 2305 379 2308 386
rect 2316 379 2319 386
rect 2363 381 2366 386
rect 2862 385 2865 392
rect 2873 385 2876 392
rect 2920 387 2923 392
rect 3017 385 3020 392
rect 3028 385 3031 392
rect 3075 387 3078 392
rect 3602 492 3604 497
rect 3621 492 3623 497
rect 3646 492 3648 497
rect 3665 492 3667 497
rect 3313 439 3316 446
rect 3324 439 3327 446
rect 3807 496 3809 501
rect 3826 496 3828 501
rect 3851 496 3853 501
rect 3870 496 3872 501
rect 5187 663 5189 668
rect 5206 663 5208 668
rect 5231 663 5233 668
rect 5250 663 5252 668
rect 3975 456 3978 463
rect 3986 456 3989 463
rect 3602 401 3605 408
rect 3613 401 3616 408
rect 3660 403 3663 408
rect 3757 401 3760 408
rect 3768 401 3771 408
rect 3815 403 3818 408
rect 3292 345 3295 352
rect 3303 345 3306 352
rect 4053 455 4056 462
rect 4064 455 4067 462
rect 4381 503 4383 508
rect 4400 503 4402 508
rect 4425 503 4427 508
rect 4444 503 4446 508
rect 4586 507 4588 512
rect 4605 507 4607 512
rect 4630 507 4632 512
rect 4649 507 4651 512
rect 4754 467 4757 474
rect 4765 467 4768 474
rect 4381 412 4384 419
rect 4392 412 4395 419
rect 4439 414 4442 419
rect 4536 412 4539 419
rect 4547 412 4550 419
rect 4594 414 4597 419
rect 4032 361 4035 368
rect 4043 361 4046 368
rect 4832 466 4835 473
rect 4843 466 4846 473
rect 5061 497 5063 502
rect 5080 497 5082 502
rect 5105 497 5107 502
rect 5124 497 5126 502
rect 5266 501 5268 506
rect 5285 501 5287 506
rect 5310 501 5312 506
rect 5329 501 5331 506
rect 5434 461 5437 468
rect 5445 461 5448 468
rect 5061 406 5064 413
rect 5072 406 5075 413
rect 5119 408 5122 413
rect 5216 406 5219 413
rect 5227 406 5230 413
rect 5274 408 5277 413
rect 4811 372 4814 379
rect 4822 372 4825 379
rect 5512 460 5515 467
rect 5523 460 5526 467
rect 5491 366 5494 373
rect 5502 366 5505 373
rect 1432 170 1435 177
rect 1443 170 1446 177
rect 1490 172 1493 177
rect 1543 172 1546 179
rect 1554 172 1557 179
rect 1601 174 1604 179
rect 1659 172 1662 179
rect 1670 172 1673 179
rect 1717 174 1720 179
rect 1779 173 1782 180
rect 1790 173 1793 180
rect 1837 175 1840 180
rect 1961 174 1964 181
rect 1972 174 1975 181
rect 2019 176 2022 181
rect 2072 176 2075 183
rect 2083 176 2086 183
rect 2130 178 2133 183
rect 2188 176 2191 183
rect 2199 176 2202 183
rect 2246 178 2249 183
rect 2308 177 2311 184
rect 2319 177 2322 184
rect 2366 179 2369 184
rect 1457 -5 1460 1
rect 1468 -5 1471 1
rect 1515 -3 1518 1
rect 1568 -5 1571 1
rect 1579 -5 1582 1
rect 1626 -3 1629 1
rect 1684 -2 1687 1
rect 1695 -2 1698 1
rect 1742 -4 1745 0
rect 1804 -1 1807 2
rect 1815 -1 1818 2
rect 1986 1 1989 4
rect 1997 1 2000 4
rect 1862 -4 1865 0
rect 2044 0 2047 4
rect 2097 3 2100 6
rect 2108 3 2111 6
rect 2155 3 2158 6
rect 2213 3 2216 6
rect 2224 3 2227 6
rect 2271 3 2274 6
rect 2333 3 2336 7
rect 2344 3 2347 7
rect 2391 3 2394 7
rect 1724 -148 1727 -141
rect 1735 -148 1738 -141
rect 1782 -146 1785 -141
rect 1842 -149 1845 -142
rect 1853 -149 1856 -142
rect 1900 -147 1903 -142
rect 1975 -149 1978 -142
rect 1986 -149 1989 -142
rect 2033 -147 2036 -142
rect 2094 -150 2097 -143
rect 2105 -150 2108 -143
rect 2152 -148 2155 -143
rect 3592 9 3595 16
rect 3603 9 3606 16
rect 3670 8 3673 15
rect 3681 8 3684 15
rect 3649 -86 3652 -79
rect 3660 -86 3663 -79
rect 3810 -118 3813 -111
rect 3821 -118 3824 -111
rect 3888 -119 3891 -112
rect 3899 -119 3902 -112
rect 3605 -267 3608 -260
rect 3616 -267 3619 -260
rect 3683 -268 3686 -261
rect 3694 -268 3697 -261
rect 4104 -153 4107 -148
rect 3867 -213 3870 -206
rect 3878 -213 3881 -206
rect 3662 -362 3665 -355
rect 3673 -362 3676 -355
rect 2837 -597 2840 -592
rect 3002 -597 3005 -592
rect 3179 -596 3182 -591
rect 3354 -597 3357 -592
rect 3752 -642 3755 -637
rect 2882 -718 2885 -711
rect 2893 -718 2896 -711
rect 2940 -716 2943 -711
rect 3053 -713 3056 -706
rect 3064 -713 3067 -706
rect 3111 -711 3114 -706
rect 3246 -717 3249 -710
rect 3257 -717 3260 -710
rect 3304 -715 3307 -710
rect 3427 -713 3430 -706
rect 3438 -713 3441 -706
rect 3485 -711 3488 -706
rect 3014 -857 3017 -850
rect 3025 -857 3028 -850
rect 3072 -855 3075 -850
rect 3018 -1055 3021 -1048
rect 3029 -1055 3032 -1048
rect 3076 -1053 3079 -1048
rect 4000 -643 4003 -638
rect 3831 -655 3833 -650
rect 3850 -655 3852 -650
rect 3875 -655 3877 -650
rect 3894 -655 3896 -650
rect 4243 -634 4246 -629
rect 4079 -656 4081 -651
rect 4098 -656 4100 -651
rect 4123 -656 4125 -651
rect 4142 -656 4144 -651
rect 4512 -629 4515 -624
rect 4322 -647 4324 -642
rect 4341 -647 4343 -642
rect 4366 -647 4368 -642
rect 4385 -647 4387 -642
rect 4591 -642 4593 -637
rect 4610 -642 4612 -637
rect 4635 -642 4637 -637
rect 4654 -642 4656 -637
rect 4085 -774 4088 -767
rect 4096 -774 4099 -767
rect 4143 -772 4146 -767
rect 4461 -786 4464 -779
rect 4472 -786 4475 -779
rect 4519 -784 4522 -779
rect 4305 -794 4308 -787
rect 4316 -794 4319 -787
rect 4363 -792 4366 -787
rect 3864 -889 3867 -882
rect 3875 -889 3878 -882
rect 3922 -887 3925 -882
rect 3877 -1075 3880 -1068
rect 3888 -1075 3891 -1068
rect 3935 -1073 3938 -1068
rect 4205 -1058 4208 -1051
rect 4216 -1058 4219 -1051
rect 4263 -1056 4266 -1051
rect 2862 -1228 2865 -1223
rect 3027 -1228 3030 -1223
rect 3204 -1227 3207 -1222
rect 3379 -1228 3382 -1223
rect 2907 -1349 2910 -1342
rect 2918 -1349 2921 -1342
rect 2965 -1347 2968 -1342
rect 3078 -1344 3081 -1337
rect 3089 -1344 3092 -1337
rect 3136 -1342 3139 -1337
rect 3271 -1348 3274 -1341
rect 3282 -1348 3285 -1341
rect 3329 -1346 3332 -1341
rect 3452 -1344 3455 -1337
rect 3463 -1344 3466 -1337
rect 3510 -1342 3513 -1337
rect 3664 -1545 3667 -1538
rect 3675 -1545 3678 -1538
rect 3742 -1546 3745 -1539
rect 3753 -1546 3756 -1539
rect 5015 -1011 5018 -1004
rect 5026 -1011 5029 -1004
rect 5073 -1009 5076 -1004
rect 5232 -1012 5235 -1005
rect 5243 -1012 5246 -1005
rect 5290 -1010 5293 -1005
rect 3721 -1640 3724 -1633
rect 3732 -1640 3735 -1633
rect 4566 -1640 4569 -1635
rect 4009 -1655 4012 -1648
rect 4020 -1655 4023 -1648
rect 3674 -1789 3677 -1782
rect 3685 -1789 3688 -1782
rect 3752 -1790 3755 -1783
rect 3763 -1790 3766 -1783
rect 4087 -1656 4090 -1649
rect 4098 -1656 4101 -1649
rect 4066 -1750 4069 -1743
rect 4077 -1750 4080 -1743
rect 3731 -1884 3734 -1877
rect 3742 -1884 3745 -1877
<< polycontact >>
rect 3035 986 3039 990
rect 3776 986 3780 990
rect 4555 986 4559 990
rect 5233 986 5237 990
rect 3035 660 3039 664
rect 3029 626 3033 630
rect 3048 626 3052 630
rect 3058 626 3062 630
rect 3776 676 3780 680
rect 3769 642 3773 646
rect 3788 642 3792 646
rect 3798 642 3802 646
rect 4555 687 4559 691
rect 4548 653 4552 657
rect 4567 653 4571 657
rect 4577 653 4581 657
rect 1297 447 1301 451
rect 1316 443 1320 447
rect 1264 424 1268 428
rect 1275 416 1279 420
rect 1271 389 1275 393
rect 1118 337 1122 341
rect 1087 314 1091 318
rect 1098 306 1102 310
rect 1145 305 1149 309
rect 2916 494 2920 498
rect 2903 460 2907 464
rect 2922 459 2926 463
rect 2932 460 2936 464
rect 1342 423 1346 427
rect 1353 415 1357 419
rect 3113 498 3117 502
rect 3108 464 3112 468
rect 3127 464 3131 468
rect 3137 464 3141 468
rect 3274 455 3278 459
rect 3234 432 3238 436
rect 3103 419 3107 423
rect 1458 385 1462 389
rect 1570 388 1574 392
rect 1685 389 1689 393
rect 1807 390 1811 394
rect 1989 391 1993 395
rect 2101 393 2105 397
rect 2217 393 2221 397
rect 2892 400 2896 404
rect 3047 400 3051 404
rect 2335 394 2339 398
rect 1316 352 1320 356
rect 1321 329 1325 333
rect 1332 321 1336 325
rect 1328 292 1332 296
rect 1140 275 1144 279
rect 1364 275 1368 280
rect 764 259 768 263
rect 1121 254 1125 258
rect 991 243 995 247
rect 1089 231 1093 235
rect 1100 223 1104 227
rect 1147 222 1151 226
rect 988 211 992 215
rect 1124 192 1128 196
rect 987 176 991 180
rect 764 150 768 154
rect 993 144 997 149
rect 989 114 993 118
rect 1118 154 1122 158
rect 1087 131 1091 135
rect 1098 123 1102 127
rect 1145 122 1149 126
rect 1128 95 1132 99
rect 989 79 994 83
rect 1119 65 1123 69
rect 1088 42 1092 46
rect 1099 34 1103 38
rect 1146 33 1150 37
rect 1124 5 1128 9
rect 1428 364 1432 368
rect 1439 356 1443 360
rect 1539 366 1543 370
rect 1486 355 1490 359
rect 1550 358 1554 362
rect 1655 366 1659 370
rect 1597 357 1601 361
rect 1666 358 1670 362
rect 1775 367 1779 371
rect 1713 357 1717 361
rect 1786 359 1790 363
rect 1957 368 1961 372
rect 1833 358 1837 362
rect 1968 360 1972 364
rect 2068 370 2072 374
rect 2015 359 2019 363
rect 2079 362 2083 366
rect 2184 370 2188 374
rect 2126 361 2130 365
rect 2195 362 2199 366
rect 2304 371 2308 375
rect 2242 361 2246 365
rect 2315 363 2319 367
rect 2861 377 2865 381
rect 2362 362 2366 366
rect 2872 369 2876 373
rect 3016 377 3020 381
rect 2919 368 2923 372
rect 3027 369 3031 373
rect 3074 368 3078 372
rect 2888 342 2892 346
rect 3245 424 3249 428
rect 3651 509 3655 513
rect 3643 476 3647 480
rect 3662 475 3666 479
rect 3672 476 3676 480
rect 3312 431 3316 435
rect 3856 514 3860 518
rect 3848 480 3852 484
rect 3867 480 3871 484
rect 3877 480 3881 484
rect 5233 681 5237 685
rect 5228 647 5232 651
rect 5247 647 5251 651
rect 5257 647 5261 651
rect 4020 471 4024 475
rect 3974 448 3978 452
rect 3849 440 3853 444
rect 3323 423 3327 427
rect 3629 416 3633 420
rect 3787 416 3791 420
rect 3601 393 3605 397
rect 3612 385 3616 389
rect 3756 393 3760 397
rect 3659 384 3663 388
rect 3767 385 3771 389
rect 3814 384 3818 388
rect 3294 363 3298 367
rect 3635 358 3639 362
rect 3791 354 3795 358
rect 3985 440 3989 444
rect 3970 413 3974 417
rect 4428 521 4432 525
rect 4422 487 4426 491
rect 4441 486 4445 490
rect 4451 487 4455 491
rect 4052 447 4056 451
rect 4633 525 4637 529
rect 4627 491 4631 495
rect 4646 491 4650 495
rect 4656 491 4660 495
rect 4789 482 4794 486
rect 4753 459 4757 463
rect 4627 449 4631 453
rect 4063 439 4067 443
rect 4409 427 4413 431
rect 4566 427 4570 431
rect 4380 404 4384 408
rect 4391 396 4395 400
rect 4535 404 4539 408
rect 4438 395 4442 399
rect 4038 379 4042 383
rect 4546 396 4550 400
rect 4593 395 4597 399
rect 4411 369 4415 373
rect 4565 365 4569 369
rect 4031 353 4035 357
rect 1461 327 1465 331
rect 1572 329 1576 333
rect 1686 329 1690 333
rect 1808 330 1812 334
rect 1990 331 1994 335
rect 2101 333 2105 337
rect 2217 333 2221 337
rect 2337 334 2341 338
rect 3046 339 3051 343
rect 3227 341 3231 345
rect 3291 337 3295 341
rect 3302 329 3306 333
rect 4042 345 4046 349
rect 4764 451 4768 455
rect 4750 424 4754 428
rect 4831 458 4835 462
rect 4842 450 4846 454
rect 5110 515 5114 519
rect 5102 481 5106 485
rect 5121 480 5125 484
rect 5131 481 5135 485
rect 5152 445 5157 450
rect 5167 445 5171 450
rect 5311 519 5315 523
rect 5307 485 5311 489
rect 5326 485 5330 489
rect 5336 485 5340 489
rect 5470 476 5474 480
rect 5433 453 5437 457
rect 5308 443 5312 447
rect 5089 421 5094 425
rect 5248 421 5253 425
rect 5060 398 5064 402
rect 4814 390 4819 394
rect 5071 390 5075 394
rect 5215 398 5219 402
rect 5118 389 5122 393
rect 5226 390 5230 394
rect 5273 389 5277 393
rect 4810 364 4814 368
rect 4821 356 4825 360
rect 5094 363 5098 367
rect 5245 362 5249 366
rect 5444 445 5448 449
rect 5435 417 5439 421
rect 5511 452 5515 456
rect 5522 444 5526 448
rect 5493 384 5497 388
rect 5490 358 5494 362
rect 4024 321 4028 325
rect 4818 327 4822 331
rect 5501 350 5505 354
rect 5501 322 5505 326
rect 1391 275 1395 280
rect 1362 82 1366 87
rect 1124 -49 1128 -45
rect 1461 185 1465 189
rect 1572 187 1576 191
rect 1688 187 1692 191
rect 1808 188 1812 192
rect 1991 189 1995 193
rect 2104 191 2108 195
rect 2219 191 2223 195
rect 2339 192 2343 196
rect 1431 162 1435 166
rect 1442 154 1446 158
rect 1542 164 1546 168
rect 1489 153 1493 157
rect 1553 156 1557 160
rect 1658 164 1662 168
rect 1600 155 1604 159
rect 1669 156 1673 160
rect 1778 165 1782 169
rect 1716 155 1720 159
rect 1789 157 1793 161
rect 1960 166 1964 170
rect 1836 156 1840 160
rect 1971 158 1975 162
rect 2071 168 2075 172
rect 2018 157 2022 161
rect 2082 160 2086 164
rect 2187 168 2191 172
rect 2129 159 2133 163
rect 2198 160 2202 164
rect 2307 169 2311 173
rect 2245 159 2249 163
rect 2318 161 2322 165
rect 2365 160 2369 164
rect 1464 125 1468 129
rect 1574 127 1578 131
rect 1691 127 1695 131
rect 1811 128 1815 132
rect 1993 129 1997 133
rect 2105 131 2109 135
rect 2220 131 2224 135
rect 2341 132 2345 136
rect 1389 82 1393 87
rect 1362 -69 1366 -64
rect 1486 8 1490 12
rect 1597 10 1601 14
rect 1712 10 1716 14
rect 1834 11 1838 15
rect 2016 12 2020 16
rect 2128 14 2132 18
rect 2245 14 2249 18
rect 2364 15 2368 19
rect 1456 -15 1460 -11
rect 1467 -23 1471 -19
rect 1567 -13 1571 -9
rect 1514 -24 1518 -20
rect 1578 -21 1582 -17
rect 1683 -13 1687 -9
rect 1625 -22 1629 -18
rect 1694 -21 1698 -17
rect 1803 -12 1807 -8
rect 1741 -22 1745 -18
rect 1814 -20 1818 -16
rect 1985 -11 1989 -7
rect 1861 -21 1865 -17
rect 1996 -19 2000 -15
rect 2096 -9 2100 -5
rect 2043 -20 2047 -16
rect 2107 -17 2111 -13
rect 2212 -9 2216 -5
rect 2154 -18 2158 -14
rect 2223 -17 2227 -13
rect 2332 -8 2336 -4
rect 2270 -18 2274 -14
rect 2343 -16 2347 -12
rect 2390 -17 2394 -13
rect 1489 -52 1493 -48
rect 1600 -50 1604 -46
rect 1715 -50 1719 -46
rect 1836 -49 1840 -45
rect 2018 -48 2022 -44
rect 2129 -46 2133 -42
rect 2245 -46 2249 -42
rect 2366 -45 2370 -41
rect 1389 -69 1393 -64
rect 1755 -133 1759 -129
rect 1871 -134 1875 -130
rect 2004 -135 2009 -131
rect 2124 -135 2128 -131
rect 1723 -156 1727 -152
rect 1734 -164 1738 -160
rect 1841 -157 1845 -153
rect 1781 -165 1785 -161
rect 1852 -165 1856 -161
rect 1974 -157 1978 -153
rect 1899 -166 1903 -162
rect 1985 -165 1989 -161
rect 2093 -158 2097 -154
rect 2032 -166 2036 -162
rect 1754 -192 1758 -188
rect 2104 -166 2108 -162
rect 2151 -167 2155 -163
rect 1873 -196 1877 -192
rect 2006 -195 2010 -191
rect 2122 -195 2126 -191
rect 2782 -215 2786 -211
rect 3631 24 3635 28
rect 3591 1 3595 5
rect 3602 -7 3606 -3
rect 3669 0 3673 4
rect 3680 -8 3684 -4
rect 3681 -35 3685 -31
rect 3654 -68 3658 -64
rect 3648 -94 3652 -90
rect 3659 -102 3663 -98
rect 3656 -131 3660 -127
rect 3839 -103 3843 -99
rect 3809 -126 3813 -122
rect 3820 -134 3824 -130
rect 3815 -162 3819 -158
rect 2827 -215 2831 -211
rect 3649 -252 3653 -248
rect 3604 -275 3608 -271
rect 3615 -283 3619 -279
rect 3610 -311 3614 -307
rect 3682 -276 3686 -272
rect 3887 -127 3891 -123
rect 3898 -135 3902 -131
rect 4108 -140 4112 -136
rect 3904 -162 3908 -158
rect 3871 -195 3875 -191
rect 3866 -221 3870 -217
rect 3877 -229 3881 -225
rect 3874 -257 3878 -253
rect 4103 -172 4107 -168
rect 4106 -207 4110 -203
rect 3693 -284 3697 -280
rect 3694 -311 3698 -307
rect 3666 -344 3670 -340
rect 3661 -370 3665 -366
rect 3672 -378 3676 -374
rect 3669 -406 3673 -402
rect 2841 -584 2845 -580
rect 2836 -616 2840 -612
rect 2821 -649 2825 -643
rect 3004 -584 3008 -580
rect 3001 -616 3005 -612
rect 3183 -583 3187 -579
rect 3178 -615 3182 -611
rect 3085 -698 3089 -694
rect 2911 -703 2915 -699
rect 3358 -584 3362 -580
rect 3353 -616 3357 -612
rect 3754 -629 3758 -625
rect 3751 -661 3755 -657
rect 3457 -698 3461 -694
rect 3737 -696 3741 -692
rect 3275 -702 3279 -698
rect 2881 -726 2885 -722
rect 2892 -734 2896 -730
rect 3052 -721 3056 -717
rect 2939 -735 2943 -731
rect 3063 -729 3067 -725
rect 3245 -725 3249 -721
rect 3110 -730 3114 -726
rect 3256 -733 3260 -729
rect 3426 -721 3430 -717
rect 3303 -734 3307 -730
rect 3437 -729 3441 -725
rect 3484 -730 3488 -726
rect 3085 -759 3089 -755
rect 3458 -759 3462 -755
rect 2913 -764 2917 -760
rect 3277 -763 3281 -759
rect 3045 -842 3049 -838
rect 3013 -865 3017 -861
rect 3024 -873 3028 -869
rect 3071 -874 3075 -870
rect 3047 -902 3051 -898
rect 3048 -1040 3052 -1036
rect 3017 -1063 3021 -1059
rect 3028 -1071 3032 -1067
rect 3075 -1072 3079 -1068
rect 3048 -1100 3052 -1096
rect 4003 -630 4007 -626
rect 3878 -637 3883 -633
rect 3872 -671 3876 -667
rect 3999 -662 4003 -658
rect 3891 -672 3895 -668
rect 3901 -671 3905 -667
rect 4006 -710 4010 -706
rect 3895 -874 3899 -870
rect 4247 -621 4251 -617
rect 4125 -638 4129 -634
rect 4242 -653 4246 -649
rect 4120 -672 4124 -668
rect 4139 -672 4143 -668
rect 4149 -672 4153 -668
rect 4514 -616 4518 -612
rect 4363 -629 4367 -625
rect 4511 -648 4515 -644
rect 4363 -663 4367 -659
rect 4382 -663 4386 -659
rect 4392 -663 4396 -659
rect 4634 -624 4638 -620
rect 4632 -658 4636 -654
rect 4651 -658 4655 -654
rect 4661 -658 4665 -654
rect 4115 -759 4119 -755
rect 4084 -782 4088 -778
rect 4095 -790 4099 -786
rect 4489 -771 4493 -767
rect 4335 -779 4339 -775
rect 4142 -791 4146 -787
rect 4304 -802 4308 -798
rect 4116 -819 4120 -815
rect 4315 -810 4319 -806
rect 4460 -794 4464 -790
rect 4362 -811 4366 -807
rect 4471 -802 4475 -798
rect 4518 -803 4522 -799
rect 4492 -831 4496 -827
rect 4336 -839 4340 -835
rect 3863 -897 3867 -893
rect 3874 -905 3878 -901
rect 3921 -906 3925 -902
rect 3895 -935 3899 -931
rect 4006 -1008 4010 -1004
rect 3905 -1060 3909 -1056
rect 4006 -1030 4010 -1026
rect 3876 -1083 3880 -1079
rect 3887 -1091 3891 -1087
rect 3934 -1092 3938 -1088
rect 3907 -1120 3911 -1116
rect 4234 -1043 4238 -1039
rect 4204 -1066 4208 -1062
rect 4215 -1074 4219 -1070
rect 4262 -1075 4266 -1071
rect 4242 -1103 4246 -1099
rect 3095 -1191 3099 -1187
rect 2864 -1215 2868 -1211
rect 2861 -1247 2865 -1243
rect 3030 -1215 3034 -1211
rect 3207 -1214 3211 -1210
rect 3382 -1215 3386 -1211
rect 3026 -1247 3030 -1243
rect 3203 -1246 3207 -1242
rect 3378 -1247 3382 -1243
rect 3107 -1329 3111 -1325
rect 2936 -1334 2940 -1330
rect 3482 -1329 3486 -1325
rect 3299 -1333 3303 -1329
rect 2906 -1357 2910 -1353
rect 2917 -1365 2921 -1361
rect 3077 -1352 3081 -1348
rect 2964 -1366 2968 -1362
rect 3088 -1360 3092 -1356
rect 3270 -1356 3274 -1352
rect 3135 -1361 3139 -1357
rect 3281 -1364 3285 -1360
rect 3451 -1352 3455 -1348
rect 3328 -1365 3332 -1361
rect 3462 -1360 3466 -1356
rect 3509 -1361 3513 -1357
rect 3110 -1390 3114 -1386
rect 3484 -1390 3488 -1386
rect 2939 -1395 2943 -1391
rect 3303 -1394 3307 -1390
rect 3705 -1530 3710 -1526
rect 3663 -1553 3667 -1549
rect 3674 -1561 3678 -1557
rect 3671 -1590 3675 -1586
rect 3741 -1554 3745 -1550
rect 3752 -1562 3756 -1558
rect 5045 -996 5049 -992
rect 5260 -997 5264 -993
rect 5014 -1019 5018 -1015
rect 5025 -1027 5029 -1023
rect 5231 -1020 5235 -1016
rect 5072 -1028 5076 -1024
rect 5242 -1028 5246 -1024
rect 5289 -1029 5293 -1025
rect 5046 -1057 5050 -1053
rect 5258 -1058 5262 -1054
rect 3757 -1589 3761 -1585
rect 3726 -1625 3731 -1621
rect 3720 -1648 3724 -1644
rect 3731 -1656 3735 -1652
rect 3729 -1685 3733 -1681
rect 4570 -1627 4574 -1623
rect 4051 -1640 4055 -1636
rect 4008 -1663 4012 -1659
rect 4019 -1671 4023 -1667
rect 4015 -1700 4019 -1696
rect 3710 -1774 3714 -1770
rect 3673 -1797 3677 -1793
rect 3684 -1805 3688 -1801
rect 3678 -1834 3682 -1830
rect 3751 -1798 3755 -1794
rect 3762 -1806 3766 -1802
rect 4086 -1664 4090 -1660
rect 4565 -1659 4569 -1655
rect 4097 -1672 4101 -1668
rect 4565 -1695 4569 -1691
rect 4094 -1701 4098 -1697
rect 4069 -1732 4073 -1728
rect 4065 -1758 4069 -1754
rect 4076 -1766 4080 -1762
rect 4073 -1795 4077 -1791
rect 3759 -1835 3763 -1831
rect 3734 -1866 3738 -1862
rect 3730 -1892 3734 -1888
rect 3741 -1900 3745 -1896
rect 3738 -1929 3742 -1925
<< ndcontact >>
rect 2983 611 2987 615
rect 2992 611 2996 615
rect 3002 611 3006 615
rect 3011 611 3015 615
rect 3027 611 3031 615
rect 3036 611 3040 615
rect 3046 611 3050 615
rect 3055 611 3059 615
rect 3723 627 3727 631
rect 3732 627 3736 631
rect 3742 627 3746 631
rect 3751 627 3755 631
rect 3767 627 3771 631
rect 3776 627 3780 631
rect 3786 627 3790 631
rect 3795 627 3799 631
rect 4502 638 4506 642
rect 4511 638 4515 642
rect 4521 638 4525 642
rect 4530 638 4534 642
rect 4546 638 4550 642
rect 4555 638 4559 642
rect 4565 638 4569 642
rect 4574 638 4578 642
rect 1259 404 1263 408
rect 1282 404 1286 408
rect 1082 294 1086 298
rect 1105 294 1109 298
rect 1138 285 1143 290
rect 1153 285 1157 290
rect 2857 445 2861 449
rect 2866 445 2870 449
rect 2876 445 2880 449
rect 2885 445 2889 449
rect 2901 445 2905 449
rect 2910 445 2914 449
rect 2920 445 2924 449
rect 2929 445 2933 449
rect 3062 449 3066 453
rect 3071 449 3075 453
rect 3081 449 3085 453
rect 3090 449 3094 453
rect 3106 449 3110 453
rect 3115 449 3119 453
rect 3125 449 3129 453
rect 3134 449 3138 453
rect 1337 403 1341 407
rect 1360 403 1364 407
rect 1316 309 1320 313
rect 1339 309 1343 313
rect 1084 211 1088 215
rect 1107 211 1111 215
rect 1140 202 1145 207
rect 1155 202 1159 207
rect 981 191 986 196
rect 996 191 1000 196
rect 982 94 987 99
rect 997 94 1001 99
rect 1082 111 1086 115
rect 1105 111 1109 115
rect 1138 102 1143 107
rect 1153 102 1157 107
rect 1083 22 1087 26
rect 1106 22 1110 26
rect 1139 13 1144 18
rect 1154 13 1158 18
rect 1423 344 1427 348
rect 1446 344 1450 348
rect 1534 346 1538 350
rect 1557 346 1561 350
rect 1650 346 1654 350
rect 1479 335 1484 340
rect 1494 335 1498 340
rect 1590 337 1595 342
rect 1605 337 1609 342
rect 1673 346 1677 350
rect 1770 347 1774 351
rect 1793 347 1797 351
rect 1952 348 1956 352
rect 1975 348 1979 352
rect 2063 350 2067 354
rect 2086 350 2090 354
rect 2179 350 2183 354
rect 1706 337 1711 342
rect 1721 337 1725 342
rect 1826 338 1831 343
rect 1841 338 1845 343
rect 2008 339 2013 344
rect 2023 339 2027 344
rect 2119 341 2124 346
rect 2134 341 2138 346
rect 2202 350 2206 354
rect 2299 351 2303 355
rect 2322 351 2326 355
rect 2856 357 2860 361
rect 2879 357 2883 361
rect 3011 357 3015 361
rect 2912 348 2917 353
rect 2927 348 2931 353
rect 3034 357 3038 361
rect 3067 348 3072 353
rect 3082 348 3086 353
rect 2235 341 2240 346
rect 2250 341 2254 346
rect 2355 342 2360 347
rect 2370 342 2374 347
rect 3229 412 3233 416
rect 3252 412 3256 416
rect 3597 461 3601 465
rect 3606 461 3610 465
rect 3616 461 3620 465
rect 3625 461 3629 465
rect 3641 461 3645 465
rect 3650 461 3654 465
rect 3660 461 3664 465
rect 3669 461 3673 465
rect 3802 465 3806 469
rect 3811 465 3815 469
rect 3821 465 3825 469
rect 3830 465 3834 469
rect 3846 465 3850 469
rect 3855 465 3859 469
rect 3865 465 3869 469
rect 3874 465 3878 469
rect 5182 632 5186 636
rect 5191 632 5195 636
rect 5201 632 5205 636
rect 5210 632 5214 636
rect 5226 632 5230 636
rect 5235 632 5239 636
rect 5245 632 5249 636
rect 5254 632 5258 636
rect 3307 411 3311 415
rect 3330 411 3334 415
rect 3596 373 3600 377
rect 3619 373 3623 377
rect 3751 373 3755 377
rect 3652 364 3657 369
rect 3667 364 3671 369
rect 3774 373 3778 377
rect 3807 364 3812 369
rect 3822 364 3826 369
rect 3969 428 3973 432
rect 3992 428 3996 432
rect 4376 472 4380 476
rect 4385 472 4389 476
rect 4395 472 4399 476
rect 4404 472 4408 476
rect 4420 472 4424 476
rect 4429 472 4433 476
rect 4439 472 4443 476
rect 4448 472 4452 476
rect 4581 476 4585 480
rect 4590 476 4594 480
rect 4600 476 4604 480
rect 4609 476 4613 480
rect 4625 476 4629 480
rect 4634 476 4638 480
rect 4644 476 4648 480
rect 4653 476 4657 480
rect 4047 427 4051 431
rect 4070 427 4074 431
rect 4375 384 4379 388
rect 4398 384 4402 388
rect 4530 384 4534 388
rect 4431 375 4436 380
rect 4446 375 4450 380
rect 4553 384 4557 388
rect 4586 375 4591 380
rect 4601 375 4605 380
rect 3286 317 3290 321
rect 3309 317 3313 321
rect 4026 333 4030 337
rect 4049 333 4053 337
rect 4748 439 4752 443
rect 4771 439 4775 443
rect 5056 466 5060 470
rect 5065 466 5069 470
rect 5075 466 5079 470
rect 5084 466 5088 470
rect 5100 466 5104 470
rect 5109 466 5113 470
rect 5119 466 5123 470
rect 5128 466 5132 470
rect 4826 438 4830 442
rect 4849 438 4853 442
rect 5261 470 5265 474
rect 5270 470 5274 474
rect 5280 470 5284 474
rect 5289 470 5293 474
rect 5305 470 5309 474
rect 5314 470 5318 474
rect 5324 470 5328 474
rect 5333 470 5337 474
rect 5055 378 5059 382
rect 5078 378 5082 382
rect 5210 378 5214 382
rect 5111 369 5116 374
rect 5126 369 5130 374
rect 5233 378 5237 382
rect 5266 369 5271 374
rect 5281 369 5285 374
rect 5428 433 5432 437
rect 5451 433 5455 437
rect 5506 432 5510 436
rect 5529 432 5533 436
rect 4805 344 4809 348
rect 4828 344 4832 348
rect 5485 338 5489 342
rect 5508 338 5512 342
rect 1426 142 1430 146
rect 1449 142 1453 146
rect 1537 144 1541 148
rect 1560 144 1564 148
rect 1653 144 1657 148
rect 1482 133 1487 138
rect 1497 133 1501 138
rect 1593 135 1598 140
rect 1608 135 1612 140
rect 1676 144 1680 148
rect 1773 145 1777 149
rect 1796 145 1800 149
rect 1955 146 1959 150
rect 1978 146 1982 150
rect 2066 148 2070 152
rect 2089 148 2093 152
rect 2182 148 2186 152
rect 1709 135 1714 140
rect 1724 135 1728 140
rect 1829 136 1834 141
rect 1844 136 1848 141
rect 2011 137 2016 142
rect 2026 137 2030 142
rect 2122 139 2127 144
rect 2137 139 2141 144
rect 2205 148 2209 152
rect 2302 149 2306 153
rect 2325 149 2329 153
rect 2238 139 2243 144
rect 2253 139 2257 144
rect 2358 140 2363 145
rect 2373 140 2377 145
rect 1451 -35 1455 -31
rect 1474 -35 1478 -31
rect 1562 -33 1566 -29
rect 1585 -33 1589 -29
rect 1678 -33 1682 -29
rect 1507 -44 1512 -39
rect 1522 -44 1526 -39
rect 1618 -42 1623 -37
rect 1633 -42 1637 -37
rect 1701 -33 1705 -29
rect 1798 -32 1802 -28
rect 1821 -32 1825 -28
rect 1980 -31 1984 -27
rect 2003 -31 2007 -27
rect 2091 -29 2095 -25
rect 2114 -29 2118 -25
rect 2207 -29 2211 -25
rect 1734 -42 1739 -37
rect 1749 -42 1753 -37
rect 1854 -41 1859 -36
rect 1869 -41 1873 -36
rect 2036 -40 2041 -35
rect 2051 -40 2055 -35
rect 2147 -38 2152 -33
rect 2162 -38 2166 -33
rect 2230 -29 2234 -25
rect 2327 -28 2331 -24
rect 2350 -28 2354 -24
rect 2263 -38 2268 -33
rect 2278 -38 2282 -33
rect 2383 -37 2388 -32
rect 2398 -37 2402 -32
rect 1718 -176 1722 -172
rect 1741 -176 1745 -172
rect 1836 -177 1840 -173
rect 1774 -185 1779 -180
rect 1789 -185 1793 -180
rect 1859 -177 1863 -173
rect 1969 -177 1973 -173
rect 1892 -186 1897 -181
rect 1907 -186 1911 -181
rect 1992 -177 1996 -173
rect 2088 -178 2092 -174
rect 2025 -186 2030 -181
rect 2040 -186 2044 -181
rect 2111 -178 2115 -174
rect 2144 -187 2149 -182
rect 2159 -187 2163 -182
rect 3586 -19 3590 -15
rect 3609 -19 3613 -15
rect 3664 -20 3668 -16
rect 3687 -20 3691 -16
rect 3643 -114 3647 -110
rect 3666 -114 3670 -110
rect 3804 -146 3808 -142
rect 3827 -146 3831 -142
rect 3599 -295 3603 -291
rect 3622 -295 3626 -291
rect 3882 -147 3886 -143
rect 3905 -147 3909 -143
rect 3861 -241 3865 -237
rect 3884 -241 3888 -237
rect 4096 -192 4101 -187
rect 4111 -192 4115 -187
rect 3677 -296 3681 -292
rect 3700 -296 3704 -292
rect 3656 -390 3660 -386
rect 3679 -390 3683 -386
rect 2829 -636 2834 -631
rect 2844 -636 2848 -631
rect 2994 -636 2999 -631
rect 3009 -636 3013 -631
rect 3171 -635 3176 -630
rect 3186 -635 3190 -630
rect 3346 -636 3351 -631
rect 3361 -636 3365 -631
rect 3744 -681 3749 -676
rect 3759 -681 3763 -676
rect 2876 -746 2880 -742
rect 2899 -746 2903 -742
rect 3047 -741 3051 -737
rect 3070 -741 3074 -737
rect 3240 -745 3244 -741
rect 3103 -750 3108 -745
rect 3118 -750 3122 -745
rect 3263 -745 3267 -741
rect 3421 -741 3425 -737
rect 3444 -741 3448 -737
rect 2932 -755 2937 -750
rect 2947 -755 2951 -750
rect 3296 -754 3301 -749
rect 3311 -754 3315 -749
rect 3477 -750 3482 -745
rect 3492 -750 3496 -745
rect 3008 -885 3012 -881
rect 3031 -885 3035 -881
rect 3064 -894 3069 -889
rect 3079 -894 3083 -889
rect 3012 -1083 3016 -1079
rect 3035 -1083 3039 -1079
rect 3068 -1092 3073 -1087
rect 3083 -1092 3087 -1087
rect 3826 -686 3830 -682
rect 3835 -686 3839 -682
rect 3845 -686 3849 -682
rect 3854 -686 3858 -682
rect 3870 -686 3874 -682
rect 3879 -686 3883 -682
rect 3889 -686 3893 -682
rect 3898 -686 3902 -682
rect 3992 -682 3997 -677
rect 4007 -682 4011 -677
rect 4074 -687 4078 -683
rect 4083 -687 4087 -683
rect 4093 -687 4097 -683
rect 4102 -687 4106 -683
rect 4118 -687 4122 -683
rect 4127 -687 4131 -683
rect 4137 -687 4141 -683
rect 4146 -687 4150 -683
rect 4235 -673 4240 -668
rect 4250 -673 4254 -668
rect 4317 -678 4321 -674
rect 4326 -678 4330 -674
rect 4336 -678 4340 -674
rect 4345 -678 4349 -674
rect 4361 -678 4365 -674
rect 4370 -678 4374 -674
rect 4380 -678 4384 -674
rect 4389 -678 4393 -674
rect 4504 -668 4509 -663
rect 4519 -668 4523 -663
rect 4586 -673 4590 -669
rect 4595 -673 4599 -669
rect 4605 -673 4609 -669
rect 4614 -673 4618 -669
rect 4630 -673 4634 -669
rect 4639 -673 4643 -669
rect 4649 -673 4653 -669
rect 4658 -673 4662 -669
rect 4079 -802 4083 -798
rect 4102 -802 4106 -798
rect 4135 -811 4140 -806
rect 4150 -811 4154 -806
rect 4299 -822 4303 -818
rect 4322 -822 4326 -818
rect 4455 -814 4459 -810
rect 4478 -814 4482 -810
rect 4511 -823 4516 -818
rect 4526 -823 4530 -818
rect 4355 -831 4360 -826
rect 4370 -831 4374 -826
rect 3858 -917 3862 -913
rect 3881 -917 3885 -913
rect 3914 -926 3919 -921
rect 3929 -926 3933 -921
rect 3871 -1103 3875 -1099
rect 3894 -1103 3898 -1099
rect 3927 -1112 3932 -1107
rect 3942 -1112 3946 -1107
rect 4199 -1086 4203 -1082
rect 4222 -1086 4226 -1082
rect 4255 -1095 4260 -1090
rect 4270 -1095 4274 -1090
rect 2854 -1267 2859 -1262
rect 2869 -1267 2873 -1262
rect 3019 -1267 3024 -1262
rect 3034 -1267 3038 -1262
rect 3196 -1266 3201 -1261
rect 3211 -1266 3215 -1261
rect 3371 -1267 3376 -1262
rect 3386 -1267 3390 -1262
rect 2901 -1377 2905 -1373
rect 2924 -1377 2928 -1373
rect 3072 -1372 3076 -1368
rect 3095 -1372 3099 -1368
rect 3265 -1376 3269 -1372
rect 3128 -1381 3133 -1376
rect 3143 -1381 3147 -1376
rect 3288 -1376 3292 -1372
rect 3446 -1372 3450 -1368
rect 3469 -1372 3473 -1368
rect 2957 -1386 2962 -1381
rect 2972 -1386 2976 -1381
rect 3321 -1385 3326 -1380
rect 3336 -1385 3340 -1380
rect 3502 -1381 3507 -1376
rect 3517 -1381 3521 -1376
rect 3658 -1573 3662 -1569
rect 3681 -1573 3685 -1569
rect 3736 -1574 3740 -1570
rect 3759 -1574 3763 -1570
rect 5009 -1039 5013 -1035
rect 5032 -1039 5036 -1035
rect 5226 -1040 5230 -1036
rect 5065 -1048 5070 -1043
rect 5080 -1048 5084 -1043
rect 5249 -1040 5253 -1036
rect 5282 -1049 5287 -1044
rect 5297 -1049 5301 -1044
rect 3715 -1668 3719 -1664
rect 3738 -1668 3742 -1664
rect 4003 -1683 4007 -1679
rect 4026 -1683 4030 -1679
rect 3668 -1817 3672 -1813
rect 3691 -1817 3695 -1813
rect 4558 -1679 4563 -1674
rect 4573 -1679 4577 -1674
rect 4081 -1684 4085 -1680
rect 4104 -1684 4108 -1680
rect 4060 -1778 4064 -1774
rect 4083 -1778 4087 -1774
rect 3746 -1818 3750 -1814
rect 3769 -1818 3773 -1814
rect 3725 -1912 3729 -1908
rect 3748 -1912 3752 -1908
<< pdcontact >>
rect 2983 642 2987 646
rect 2992 642 2996 646
rect 3002 642 3006 646
rect 3011 642 3015 646
rect 3027 642 3031 646
rect 3036 642 3040 646
rect 3046 642 3050 646
rect 3055 642 3059 646
rect 3723 658 3727 662
rect 3732 658 3736 662
rect 3742 658 3746 662
rect 3751 658 3755 662
rect 3767 658 3771 662
rect 3776 658 3780 662
rect 3786 658 3790 662
rect 3795 658 3799 662
rect 4502 669 4506 673
rect 4511 669 4515 673
rect 4521 669 4525 673
rect 4530 669 4534 673
rect 4546 669 4550 673
rect 4555 669 4559 673
rect 4565 669 4569 673
rect 4574 669 4578 673
rect 1258 435 1262 439
rect 1271 435 1275 439
rect 1282 435 1286 439
rect 1081 325 1085 329
rect 1094 325 1098 329
rect 1105 325 1109 329
rect 1138 324 1142 329
rect 1153 324 1157 329
rect 1336 434 1340 438
rect 1349 434 1353 438
rect 1360 434 1364 438
rect 2857 476 2861 480
rect 2866 476 2870 480
rect 2876 476 2880 480
rect 2885 476 2889 480
rect 2901 476 2905 480
rect 2910 476 2914 480
rect 2920 476 2924 480
rect 2929 476 2933 480
rect 3062 480 3066 484
rect 3071 480 3075 484
rect 3081 480 3085 484
rect 3090 480 3094 484
rect 3106 480 3110 484
rect 3115 480 3119 484
rect 3125 480 3129 484
rect 3134 480 3138 484
rect 3228 443 3232 447
rect 3241 443 3245 447
rect 3252 443 3256 447
rect 2855 388 2859 392
rect 1315 340 1319 344
rect 1328 340 1332 344
rect 1339 340 1343 344
rect 1083 242 1087 246
rect 1096 242 1100 246
rect 1107 242 1111 246
rect 1140 241 1144 246
rect 1155 241 1159 246
rect 981 230 985 235
rect 996 230 1000 235
rect 982 133 986 138
rect 997 133 1001 138
rect 1081 142 1085 146
rect 1094 142 1098 146
rect 1105 142 1109 146
rect 1138 141 1142 146
rect 1153 141 1157 146
rect 1082 53 1086 57
rect 1095 53 1099 57
rect 1106 53 1110 57
rect 1139 52 1143 57
rect 1154 52 1158 57
rect 1422 375 1426 379
rect 1435 375 1439 379
rect 1446 375 1450 379
rect 1479 374 1483 379
rect 1494 374 1498 379
rect 1533 377 1537 381
rect 1546 377 1550 381
rect 1557 377 1561 381
rect 1590 376 1594 381
rect 1605 376 1609 381
rect 1649 377 1653 381
rect 1662 377 1666 381
rect 1673 377 1677 381
rect 1706 376 1710 381
rect 1721 376 1725 381
rect 1769 378 1773 382
rect 1782 378 1786 382
rect 1793 378 1797 382
rect 1826 377 1830 382
rect 1841 377 1845 382
rect 1951 379 1955 383
rect 1964 379 1968 383
rect 1975 379 1979 383
rect 2008 378 2012 383
rect 2023 378 2027 383
rect 2062 381 2066 385
rect 2075 381 2079 385
rect 2086 381 2090 385
rect 2119 380 2123 385
rect 2134 380 2138 385
rect 2178 381 2182 385
rect 2191 381 2195 385
rect 2202 381 2206 385
rect 2235 380 2239 385
rect 2250 380 2254 385
rect 2298 382 2302 386
rect 2311 382 2315 386
rect 2322 382 2326 386
rect 2355 381 2359 386
rect 2370 381 2374 386
rect 2868 388 2872 392
rect 2879 388 2883 392
rect 2912 387 2916 392
rect 2927 387 2931 392
rect 3010 388 3014 392
rect 3023 388 3027 392
rect 3034 388 3038 392
rect 3067 387 3071 392
rect 3082 387 3086 392
rect 3597 492 3601 496
rect 3606 492 3610 496
rect 3616 492 3620 496
rect 3625 492 3629 496
rect 3641 492 3645 496
rect 3650 492 3654 496
rect 3660 492 3664 496
rect 3669 492 3673 496
rect 3306 442 3310 446
rect 3319 442 3323 446
rect 3330 442 3334 446
rect 3802 496 3806 500
rect 3811 496 3815 500
rect 3821 496 3825 500
rect 3830 496 3834 500
rect 3846 496 3850 500
rect 3855 496 3859 500
rect 3865 496 3869 500
rect 3874 496 3878 500
rect 5182 663 5186 667
rect 5191 663 5195 667
rect 5201 663 5205 667
rect 5210 663 5214 667
rect 5226 663 5230 667
rect 5235 663 5239 667
rect 5245 663 5249 667
rect 5254 663 5258 667
rect 3968 459 3972 463
rect 3981 459 3985 463
rect 3992 459 3996 463
rect 3595 404 3599 408
rect 3608 404 3612 408
rect 3619 404 3623 408
rect 3652 403 3656 408
rect 3667 403 3671 408
rect 3750 404 3754 408
rect 3763 404 3767 408
rect 3774 404 3778 408
rect 3807 403 3811 408
rect 3822 403 3826 408
rect 3285 348 3289 352
rect 3298 348 3302 352
rect 3309 348 3313 352
rect 4046 458 4050 462
rect 4059 458 4063 462
rect 4070 458 4074 462
rect 4376 503 4380 507
rect 4385 503 4389 507
rect 4395 503 4399 507
rect 4404 503 4408 507
rect 4420 503 4424 507
rect 4429 503 4433 507
rect 4439 503 4443 507
rect 4448 503 4452 507
rect 4581 507 4585 511
rect 4590 507 4594 511
rect 4600 507 4604 511
rect 4609 507 4613 511
rect 4625 507 4629 511
rect 4634 507 4638 511
rect 4644 507 4648 511
rect 4653 507 4657 511
rect 4747 470 4751 474
rect 4760 470 4764 474
rect 4771 470 4775 474
rect 4374 415 4378 419
rect 4387 415 4391 419
rect 4398 415 4402 419
rect 4431 414 4435 419
rect 4446 414 4450 419
rect 4529 415 4533 419
rect 4542 415 4546 419
rect 4553 415 4557 419
rect 4586 414 4590 419
rect 4601 414 4605 419
rect 4025 364 4029 368
rect 4038 364 4042 368
rect 4049 364 4053 368
rect 4825 469 4829 473
rect 4838 469 4842 473
rect 4849 469 4853 473
rect 5056 497 5060 501
rect 5065 497 5069 501
rect 5075 497 5079 501
rect 5084 497 5088 501
rect 5100 497 5104 501
rect 5109 497 5113 501
rect 5119 497 5123 501
rect 5128 497 5132 501
rect 5261 501 5265 505
rect 5270 501 5274 505
rect 5280 501 5284 505
rect 5289 501 5293 505
rect 5305 501 5309 505
rect 5314 501 5318 505
rect 5324 501 5328 505
rect 5333 501 5337 505
rect 5427 464 5431 468
rect 5440 464 5444 468
rect 5451 464 5455 468
rect 5054 409 5058 413
rect 5067 409 5071 413
rect 5078 409 5082 413
rect 5111 408 5115 413
rect 5126 408 5130 413
rect 5209 409 5213 413
rect 5222 409 5226 413
rect 5233 409 5237 413
rect 5266 408 5270 413
rect 5281 408 5285 413
rect 4804 375 4808 379
rect 4817 375 4821 379
rect 4828 375 4832 379
rect 5505 463 5509 467
rect 5518 463 5522 467
rect 5529 463 5533 467
rect 5484 369 5488 373
rect 5497 369 5501 373
rect 5508 369 5512 373
rect 1425 173 1429 177
rect 1438 173 1442 177
rect 1449 173 1453 177
rect 1482 172 1486 177
rect 1497 172 1501 177
rect 1536 175 1540 179
rect 1549 175 1553 179
rect 1560 175 1564 179
rect 1593 174 1597 179
rect 1608 174 1612 179
rect 1652 175 1656 179
rect 1665 175 1669 179
rect 1676 175 1680 179
rect 1709 174 1713 179
rect 1724 174 1728 179
rect 1772 176 1776 180
rect 1785 176 1789 180
rect 1796 176 1800 180
rect 1829 175 1833 180
rect 1844 175 1848 180
rect 1954 177 1958 181
rect 1967 177 1971 181
rect 1978 177 1982 181
rect 2011 176 2015 181
rect 2026 176 2030 181
rect 2065 179 2069 183
rect 2078 179 2082 183
rect 2089 179 2093 183
rect 2122 178 2126 183
rect 2137 178 2141 183
rect 2181 179 2185 183
rect 2194 179 2198 183
rect 2205 179 2209 183
rect 2238 178 2242 183
rect 2253 178 2257 183
rect 2301 180 2305 184
rect 2314 180 2318 184
rect 2325 180 2329 184
rect 2358 179 2362 184
rect 2373 179 2377 184
rect 1450 -2 1454 2
rect 1463 -2 1467 2
rect 1474 -2 1478 2
rect 1507 -3 1511 1
rect 1522 -3 1526 1
rect 1561 -2 1565 2
rect 1574 -2 1578 2
rect 1585 -2 1589 2
rect 1618 -3 1622 1
rect 1633 -3 1637 1
rect 1677 -2 1681 2
rect 1690 -2 1694 2
rect 1701 -2 1705 2
rect 1734 -4 1738 0
rect 1749 -4 1753 0
rect 1797 -1 1801 3
rect 1810 -1 1814 3
rect 1821 -1 1825 3
rect 1979 1 1983 5
rect 1992 1 1996 5
rect 2003 1 2007 5
rect 1854 -4 1858 0
rect 1869 -4 1873 0
rect 2036 0 2040 4
rect 2051 0 2055 4
rect 2090 3 2094 7
rect 2103 3 2107 7
rect 2114 3 2118 7
rect 2147 3 2151 7
rect 2162 3 2166 7
rect 2206 3 2210 7
rect 2219 3 2223 7
rect 2230 3 2234 7
rect 2263 2 2267 6
rect 2278 3 2282 7
rect 2326 3 2330 7
rect 2339 3 2343 7
rect 2350 3 2354 7
rect 2383 3 2387 7
rect 2398 3 2402 7
rect 1717 -145 1721 -141
rect 1730 -145 1734 -141
rect 1741 -145 1745 -141
rect 1774 -146 1778 -141
rect 1789 -146 1793 -141
rect 1835 -146 1839 -142
rect 1848 -146 1852 -142
rect 1859 -146 1863 -142
rect 1892 -147 1896 -142
rect 1907 -147 1911 -142
rect 1968 -146 1972 -142
rect 1981 -146 1985 -142
rect 1992 -146 1996 -142
rect 2025 -147 2029 -142
rect 2040 -147 2044 -142
rect 2087 -147 2091 -143
rect 2100 -147 2104 -143
rect 2111 -147 2115 -143
rect 2144 -148 2148 -143
rect 2159 -148 2163 -143
rect 3585 12 3589 16
rect 3598 12 3602 16
rect 3609 12 3613 16
rect 3663 11 3667 15
rect 3676 11 3680 15
rect 3687 11 3691 15
rect 3642 -83 3646 -79
rect 3655 -83 3659 -79
rect 3666 -83 3670 -79
rect 3803 -115 3807 -111
rect 3816 -115 3820 -111
rect 3827 -115 3831 -111
rect 3881 -116 3885 -112
rect 3894 -116 3898 -112
rect 3905 -116 3909 -112
rect 3598 -264 3602 -260
rect 3611 -264 3615 -260
rect 3622 -264 3626 -260
rect 3676 -265 3680 -261
rect 3689 -265 3693 -261
rect 3700 -265 3704 -261
rect 4096 -153 4100 -148
rect 4111 -153 4115 -148
rect 3860 -210 3864 -206
rect 3873 -210 3877 -206
rect 3884 -210 3888 -206
rect 3655 -359 3659 -355
rect 3668 -359 3672 -355
rect 3679 -359 3683 -355
rect 2829 -597 2833 -592
rect 2844 -597 2848 -592
rect 2994 -597 2998 -592
rect 3009 -597 3013 -592
rect 3171 -596 3175 -591
rect 3186 -596 3190 -591
rect 3346 -597 3350 -592
rect 3361 -597 3365 -592
rect 3744 -642 3748 -637
rect 3759 -642 3763 -637
rect 3046 -710 3050 -706
rect 2875 -715 2879 -711
rect 2888 -715 2892 -711
rect 2899 -715 2903 -711
rect 2932 -716 2936 -711
rect 2947 -716 2951 -711
rect 3059 -710 3063 -706
rect 3070 -710 3074 -706
rect 3103 -711 3107 -706
rect 3118 -711 3122 -706
rect 3420 -710 3424 -706
rect 3239 -714 3243 -710
rect 3252 -714 3256 -710
rect 3263 -714 3267 -710
rect 3296 -715 3300 -710
rect 3311 -715 3315 -710
rect 3433 -710 3437 -706
rect 3444 -710 3448 -706
rect 3477 -711 3481 -706
rect 3492 -711 3496 -706
rect 3007 -854 3011 -850
rect 3020 -854 3024 -850
rect 3031 -854 3035 -850
rect 3064 -855 3068 -850
rect 3079 -855 3083 -850
rect 3011 -1052 3015 -1048
rect 3024 -1052 3028 -1048
rect 3035 -1052 3039 -1048
rect 3068 -1053 3072 -1048
rect 3083 -1053 3087 -1048
rect 3992 -643 3996 -638
rect 4007 -643 4011 -638
rect 3826 -655 3830 -651
rect 3835 -655 3839 -651
rect 3845 -655 3849 -651
rect 3854 -655 3858 -651
rect 3870 -655 3874 -651
rect 3879 -655 3883 -651
rect 3889 -655 3893 -651
rect 3898 -655 3902 -651
rect 4235 -634 4239 -629
rect 4250 -634 4254 -629
rect 4074 -656 4078 -652
rect 4083 -656 4087 -652
rect 4093 -656 4097 -652
rect 4102 -656 4106 -652
rect 4118 -656 4122 -652
rect 4127 -656 4131 -652
rect 4137 -656 4141 -652
rect 4146 -656 4150 -652
rect 4504 -629 4508 -624
rect 4519 -629 4523 -624
rect 4317 -647 4321 -643
rect 4326 -647 4330 -643
rect 4336 -647 4340 -643
rect 4345 -647 4349 -643
rect 4361 -647 4365 -643
rect 4370 -647 4374 -643
rect 4380 -647 4384 -643
rect 4389 -647 4393 -643
rect 4586 -642 4590 -638
rect 4595 -642 4599 -638
rect 4605 -642 4609 -638
rect 4614 -642 4618 -638
rect 4630 -642 4634 -638
rect 4639 -642 4643 -638
rect 4649 -642 4653 -638
rect 4658 -642 4662 -638
rect 4078 -771 4082 -767
rect 4091 -771 4095 -767
rect 4102 -771 4106 -767
rect 4135 -772 4139 -767
rect 4150 -772 4154 -767
rect 4454 -783 4458 -779
rect 4467 -783 4471 -779
rect 4478 -783 4482 -779
rect 4511 -784 4515 -779
rect 4526 -784 4530 -779
rect 4298 -791 4302 -787
rect 4311 -791 4315 -787
rect 4322 -791 4326 -787
rect 4355 -792 4359 -787
rect 4370 -792 4374 -787
rect 3857 -886 3861 -882
rect 3870 -886 3874 -882
rect 3881 -886 3885 -882
rect 3914 -887 3918 -882
rect 3929 -887 3933 -882
rect 3870 -1072 3874 -1068
rect 3883 -1072 3887 -1068
rect 3894 -1072 3898 -1068
rect 3927 -1073 3931 -1068
rect 3942 -1073 3946 -1068
rect 4198 -1055 4202 -1051
rect 4211 -1055 4215 -1051
rect 4222 -1055 4226 -1051
rect 4255 -1056 4259 -1051
rect 4270 -1056 4274 -1051
rect 2854 -1228 2858 -1223
rect 2869 -1228 2873 -1223
rect 3019 -1228 3023 -1223
rect 3034 -1228 3038 -1223
rect 3196 -1227 3200 -1222
rect 3211 -1227 3215 -1222
rect 3371 -1228 3375 -1223
rect 3386 -1228 3390 -1223
rect 3071 -1341 3075 -1337
rect 2900 -1346 2904 -1342
rect 2913 -1346 2917 -1342
rect 2924 -1346 2928 -1342
rect 2957 -1347 2961 -1342
rect 2972 -1347 2976 -1342
rect 3084 -1341 3088 -1337
rect 3095 -1341 3099 -1337
rect 3128 -1342 3132 -1337
rect 3143 -1342 3147 -1337
rect 3445 -1341 3449 -1337
rect 3264 -1345 3268 -1341
rect 3277 -1345 3281 -1341
rect 3288 -1345 3292 -1341
rect 3321 -1346 3325 -1341
rect 3336 -1346 3340 -1341
rect 3458 -1341 3462 -1337
rect 3469 -1341 3473 -1337
rect 3502 -1342 3506 -1337
rect 3517 -1342 3521 -1337
rect 3657 -1542 3661 -1538
rect 3670 -1542 3674 -1538
rect 3681 -1542 3685 -1538
rect 3735 -1543 3739 -1539
rect 3748 -1543 3752 -1539
rect 3759 -1543 3763 -1539
rect 5008 -1008 5012 -1004
rect 5021 -1008 5025 -1004
rect 5032 -1008 5036 -1004
rect 5065 -1009 5069 -1004
rect 5080 -1009 5084 -1004
rect 5225 -1009 5229 -1005
rect 5238 -1009 5242 -1005
rect 5249 -1009 5253 -1005
rect 5282 -1010 5286 -1005
rect 5297 -1010 5301 -1005
rect 3714 -1637 3718 -1633
rect 3727 -1637 3731 -1633
rect 3738 -1637 3742 -1633
rect 4558 -1640 4562 -1635
rect 4573 -1640 4577 -1635
rect 4002 -1652 4006 -1648
rect 4015 -1652 4019 -1648
rect 4026 -1652 4030 -1648
rect 3667 -1786 3671 -1782
rect 3680 -1786 3684 -1782
rect 3691 -1786 3695 -1782
rect 3745 -1787 3749 -1783
rect 3758 -1787 3762 -1783
rect 3769 -1787 3773 -1783
rect 4080 -1653 4084 -1649
rect 4093 -1653 4097 -1649
rect 4104 -1653 4108 -1649
rect 4059 -1747 4063 -1743
rect 4072 -1747 4076 -1743
rect 4083 -1747 4087 -1743
rect 3724 -1881 3728 -1877
rect 3737 -1881 3741 -1877
rect 3748 -1881 3752 -1877
<< m2contact >>
rect 5239 833 5243 837
rect 4100 771 4104 775
rect 3360 755 3364 759
rect 964 211 968 215
rect 1328 423 1332 427
rect 1281 389 1285 393
rect 1348 387 1352 391
rect 1417 356 1421 360
rect 1528 358 1532 362
rect 1077 231 1081 235
rect 1044 131 1049 135
rect 1160 222 1165 226
rect 1644 358 1648 362
rect 1764 359 1769 363
rect 1946 360 1950 364
rect 2026 359 2030 363
rect 2057 362 2061 366
rect 2137 362 2141 366
rect 2173 362 2177 366
rect 2252 360 2256 364
rect 2296 363 2300 367
rect 2996 663 3000 667
rect 3043 626 3047 630
rect 2885 497 2889 501
rect 2918 453 2922 457
rect 3092 508 3096 512
rect 3122 457 3126 461
rect 2849 369 2854 373
rect 3004 377 3009 381
rect 3004 369 3008 373
rect 3088 369 3092 373
rect 3300 431 3304 435
rect 3239 396 3243 400
rect 3318 396 3322 400
rect 3753 688 3757 693
rect 3736 679 3740 683
rect 3783 642 3787 646
rect 3625 513 3629 517
rect 3658 469 3662 473
rect 3832 524 3836 528
rect 3862 473 3866 477
rect 3552 393 3556 397
rect 3589 385 3594 389
rect 3744 393 3749 397
rect 3744 385 3748 389
rect 3828 385 3832 389
rect 4040 447 4044 451
rect 3986 412 3990 416
rect 4045 412 4049 416
rect 4534 698 4538 703
rect 4515 690 4519 694
rect 4562 653 4566 657
rect 4404 524 4408 528
rect 4437 480 4441 484
rect 4611 535 4615 539
rect 4641 484 4645 488
rect 4330 404 4335 408
rect 4368 396 4373 400
rect 4523 404 4528 408
rect 4523 396 4527 400
rect 4607 396 4611 400
rect 4819 458 4823 462
rect 4758 423 4762 427
rect 4837 422 4841 426
rect 5084 518 5088 522
rect 5117 474 5121 478
rect 3550 251 3554 255
rect 4328 238 4332 243
rect 5048 390 5053 394
rect 5211 693 5215 697
rect 5195 684 5199 688
rect 5240 690 5244 695
rect 5242 647 5246 651
rect 5291 529 5295 533
rect 5321 485 5325 489
rect 5203 398 5208 402
rect 5287 390 5291 394
rect 5499 452 5503 456
rect 5442 417 5446 421
rect 5517 416 5521 420
rect 5520 352 5525 356
rect 1076 131 1081 135
rect 1420 154 1424 158
rect 1531 156 1535 160
rect 1078 42 1082 46
rect 1647 156 1651 160
rect 1767 157 1771 161
rect 1949 158 1953 162
rect 2033 157 2037 161
rect 2060 160 2064 164
rect 2143 158 2147 163
rect 2176 160 2180 164
rect 2260 159 2265 163
rect 2296 161 2300 165
rect 2380 160 2384 164
rect 1445 -23 1449 -19
rect 1556 -21 1560 -17
rect 1672 -21 1676 -17
rect 1792 -20 1796 -16
rect 1974 -19 1978 -15
rect 1712 -164 1716 -160
rect 1819 -165 1823 -161
rect 2085 -17 2089 -13
rect 2201 -17 2205 -13
rect 2323 -16 2327 -12
rect 2182 -54 2186 -50
rect 2062 -65 2066 -61
rect 1963 -165 1967 -161
rect 2287 -208 2291 -204
rect 3575 1 3581 5
rect 3654 -1 3661 4
rect 3672 -100 3676 -96
rect 3588 -275 3594 -271
rect 3667 -277 3674 -272
rect 3872 -128 3879 -123
rect 2762 -534 2769 -530
rect 2764 -555 2768 -551
rect 2764 -571 2768 -567
rect 2764 -616 2769 -611
rect 2707 -669 2712 -665
rect 2806 -669 2810 -665
rect 2708 -682 2713 -678
rect 2792 -682 2796 -678
rect 2710 -696 2715 -692
rect 2773 -696 2777 -692
rect 2713 -735 2717 -731
rect 2758 -735 2762 -731
rect 2830 -616 2835 -611
rect 2834 -652 2838 -648
rect 2842 -736 2846 -732
rect 2996 -616 3000 -612
rect 3171 -615 3176 -611
rect 3001 -652 3006 -648
rect 2870 -734 2874 -730
rect 3178 -651 3183 -647
rect 3021 -731 3025 -727
rect 3041 -729 3045 -725
rect 3348 -616 3352 -612
rect 3353 -652 3357 -648
rect 2956 -821 2960 -817
rect 3123 -729 3127 -725
rect 3210 -735 3214 -731
rect 3234 -733 3239 -729
rect 3415 -729 3419 -725
rect 3497 -729 3501 -725
rect 3324 -734 3329 -730
rect 4132 -582 4136 -578
rect 4375 -593 4379 -588
rect 4645 -595 4649 -591
rect 3862 -626 3866 -622
rect 4346 -619 4350 -614
rect 4618 -613 4622 -609
rect 3746 -661 3750 -657
rect 3751 -697 3756 -693
rect 2984 -821 2988 -817
rect 3838 -634 3842 -630
rect 4105 -627 4109 -623
rect 3994 -662 3998 -658
rect 4010 -662 4015 -658
rect 3886 -672 3890 -668
rect 4086 -635 4090 -631
rect 4237 -653 4241 -649
rect 4134 -672 4138 -668
rect 3875 -693 3879 -689
rect 4244 -689 4248 -685
rect 4329 -626 4333 -622
rect 4506 -648 4510 -644
rect 4377 -663 4381 -659
rect 4598 -621 4602 -617
rect 4646 -658 4650 -654
rect 4369 -685 4373 -681
rect 4070 -783 4074 -779
rect 3085 -873 3089 -869
rect 3849 -898 3853 -894
rect 2978 -1169 2983 -1165
rect 2978 -1184 2983 -1180
rect 2858 -1282 2862 -1278
rect 2982 -1247 2986 -1243
rect 2896 -1365 2900 -1361
rect 3089 -1071 3093 -1067
rect 3934 -905 3938 -901
rect 4290 -803 4294 -799
rect 4376 -810 4380 -806
rect 3015 -1169 3021 -1165
rect 3013 -1184 3020 -1180
rect 3021 -1247 3025 -1243
rect 3025 -1283 3029 -1279
rect 3203 -1282 3207 -1278
rect 3094 -1290 3098 -1286
rect 3066 -1360 3070 -1356
rect 3378 -1283 3382 -1279
rect 3260 -1364 3264 -1360
rect 3439 -1360 3445 -1356
rect 3523 -1360 3527 -1356
rect 3948 -1091 3952 -1087
rect 4277 -1075 4285 -1069
rect 3647 -1553 3653 -1549
rect 3726 -1555 3733 -1550
rect 3744 -1654 3748 -1650
rect 3657 -1797 3663 -1793
rect 3736 -1799 3743 -1794
rect 4071 -1665 4078 -1660
<< m3contact >>
rect 2050 362 2054 366
rect 2161 362 2166 366
rect 2283 363 2288 367
rect 2050 160 2054 164
rect 2161 160 2166 164
rect 2283 161 2288 165
rect 2074 -17 2078 -13
rect 2194 -17 2198 -13
rect 2315 -16 2320 -12
rect 3306 -534 3310 -530
rect 3145 -555 3149 -551
rect 2958 -571 2962 -567
rect 2775 -618 2779 -613
rect 2974 -619 2978 -614
rect 3154 -618 3158 -613
rect 3332 -619 3336 -614
rect 3860 -537 3866 -530
rect 4103 -557 4109 -550
rect 4345 -574 4351 -567
rect 4618 -566 4623 -561
rect 3036 -1364 3041 -1358
rect 3405 -1361 3410 -1355
rect 3227 -1370 3232 -1364
rect 2867 -1382 2872 -1376
<< nsubstratencontact >>
rect 1141 335 1145 339
rect 1482 385 1486 389
rect 1593 387 1597 391
rect 1709 387 1713 391
rect 1829 388 1833 392
rect 2011 389 2015 393
rect 2122 391 2126 395
rect 2915 398 2919 402
rect 3070 398 3074 402
rect 2238 391 2242 395
rect 2358 392 2362 396
rect 1143 252 1147 256
rect 984 241 988 245
rect 985 144 989 148
rect 1141 152 1145 156
rect 1142 63 1146 67
rect 3655 414 3659 418
rect 3810 414 3814 418
rect 4434 425 4438 429
rect 4589 425 4593 429
rect 5114 419 5118 423
rect 5269 419 5273 423
rect 1485 183 1489 187
rect 1596 185 1600 189
rect 1712 185 1716 189
rect 1832 186 1836 190
rect 2014 187 2018 191
rect 2125 189 2129 193
rect 2241 189 2245 193
rect 2361 190 2365 194
rect 1510 6 1514 10
rect 1621 8 1625 12
rect 1737 8 1741 12
rect 1857 9 1861 13
rect 2039 10 2043 14
rect 2150 12 2154 16
rect 2266 12 2270 16
rect 2386 13 2390 17
rect 1777 -135 1781 -131
rect 1895 -136 1899 -132
rect 2028 -136 2032 -132
rect 2147 -137 2151 -133
rect 4099 -142 4103 -138
rect 2832 -586 2836 -582
rect 2997 -586 3001 -582
rect 3174 -585 3178 -581
rect 3106 -700 3110 -696
rect 3349 -586 3353 -582
rect 3747 -631 3751 -627
rect 2935 -705 2939 -701
rect 3480 -700 3484 -696
rect 3299 -704 3303 -700
rect 3067 -844 3071 -840
rect 3071 -1042 3075 -1038
rect 3995 -632 3999 -628
rect 4238 -623 4242 -619
rect 4507 -618 4511 -614
rect 4138 -761 4142 -757
rect 4514 -773 4518 -769
rect 4358 -781 4362 -777
rect 3917 -876 3921 -872
rect 3930 -1062 3934 -1058
rect 4258 -1045 4262 -1041
rect 2857 -1217 2861 -1213
rect 3022 -1217 3026 -1213
rect 3199 -1216 3203 -1212
rect 3374 -1217 3378 -1213
rect 3131 -1331 3135 -1327
rect 2960 -1336 2964 -1332
rect 3505 -1331 3509 -1327
rect 3324 -1335 3328 -1331
rect 5068 -998 5072 -994
rect 5285 -999 5289 -995
rect 4561 -1629 4565 -1625
<< labels >>
rlabel metal1 1155 308 1155 308 1 D0
rlabel metal1 1157 224 1157 224 1 D1
rlabel metal1 1156 124 1156 124 1 D2
rlabel metal1 1156 33 1156 33 1 D3
rlabel metal1 978 213 978 213 1 S0
rlabel metal1 980 117 980 117 1 S1
rlabel metal1 1951 362 1951 362 1 B0
rlabel metal1 2026 360 2026 360 1 b1_f_0
rlabel metal1 2062 363 2062 363 1 B1
rlabel metal1 2137 363 2137 363 1 b1_f_1
rlabel metal1 2178 363 2178 363 1 B2
rlabel metal1 2252 362 2252 362 1 b1_f_2
rlabel m2contact 2299 365 2299 365 1 B3
rlabel metal1 2372 363 2372 363 1 b1_f_3
rlabel metal1 1844 358 1844 358 1 a1_f_3
rlabel metal1 1724 359 1724 359 1 a1_f_2
rlabel metal1 1496 357 1496 357 1 a1_f_0
rlabel metal1 1769 362 1769 362 1 A3
rlabel metal1 1650 359 1650 359 1 A2
rlabel metal1 1534 360 1534 360 1 A1
rlabel metal1 1421 358 1421 358 1 A0
rlabel metal1 1500 155 1500 155 1 a2_f_0
rlabel metal1 1611 157 1611 157 1 a2_f_1
rlabel metal1 1726 157 1726 157 1 a2_f_2
rlabel metal1 1846 156 1846 156 1 a2_f_3
rlabel metal1 1525 -21 1525 -21 1 a3_f_0
rlabel metal1 1635 -19 1635 -19 1 a3_f_1
rlabel metal1 1752 -19 1752 -19 1 a3_f_2
rlabel metal1 1871 -19 1871 -19 1 a3_f_3
rlabel metal1 1409 395 1409 395 1 deff
rlabel metal1 2028 159 2028 159 1 b2_f_0
rlabel metal1 2139 162 2139 162 1 b2_f_1
rlabel metal1 2255 162 2255 162 1 b2_f_2
rlabel metal1 2375 162 2375 162 1 b2_f_3
rlabel metal1 2053 -19 2053 -19 1 b3_f_0
rlabel metal1 2164 -16 2164 -16 1 b3_f_1
rlabel metal1 2280 -15 2280 -15 1 b3_f_2
rlabel metal1 2400 -16 2400 -16 1 b3_f_3
rlabel m2contact 5521 354 5521 354 1 C1
rlabel metal1 3324 333 3324 333 1 carry
rlabel metal1 4062 350 4062 350 1 C3
rlabel metal1 4841 361 4841 361 1 C2
rlabel metal1 3078 503 3078 503 1 sum_3
rlabel metal1 3818 519 3818 519 1 sum_2
rlabel metal1 4596 529 4596 529 1 sum_1
rlabel metal1 5275 524 5275 524 1 sum_0
rlabel metal1 1794 -162 1794 -162 1 a4_0
rlabel metal1 1911 -163 1911 -163 1 a4_1
rlabel metal1 2044 -163 2044 -163 1 a4_2
rlabel metal1 2164 -164 2164 -164 1 a4_3
rlabel metal1 2846 -614 2846 -614 1 na0
rlabel metal1 3011 -614 3011 -614 1 na1
rlabel metal1 2951 -732 2951 -732 1 w7
rlabel metal1 3121 -728 3121 -728 1 w5
rlabel metal1 3363 -615 3363 -615 1 na3
rlabel metal1 3497 -728 3497 -728 1 w1
rlabel metal1 3314 -731 3314 -731 1 w3
rlabel metal1 3188 -614 3188 -614 1 na2
rlabel metal1 3762 -661 3762 -661 1 x3
rlabel metal1 4009 -661 4009 -661 1 x2
rlabel metal1 4252 -653 4252 -653 1 x1
rlabel metal1 4522 -648 4522 -648 1 x0
rlabel metal1 2872 -1244 2872 -1244 1 nb0
rlabel metal1 3042 -1244 3042 -1244 1 nb1
rlabel metal1 3217 -1243 3217 -1243 1 nb2
rlabel metal1 3392 -1245 3392 -1245 1 nb3
rlabel metal1 2977 -1363 2977 -1363 1 w8
rlabel metal1 3341 -1362 3341 -1362 1 w4
rlabel metal1 3521 -1358 3521 -1358 1 w2
rlabel metal1 3933 -903 3933 -903 1 t1
rlabel metal1 3947 -1089 3947 -1089 1 t2
rlabel metal1 4153 -788 4153 -788 1 o1
rlabel metal1 4374 -808 4374 -808 1 t3
rlabel metal1 3148 -1358 3148 -1358 1 w6
rlabel metal1 4274 -1073 4274 -1073 1 t4
rlabel metal1 4531 -801 4531 -801 1 o2
rlabel metal1 3083 -872 3083 -872 1 t5
rlabel metal1 3089 -1069 3089 -1069 1 t6
rlabel metal1 3685 -375 3685 -375 1 l1
rlabel metal1 3671 -98 3671 -98 1 l2
rlabel metal1 3742 -1652 3742 -1652 1 g1
rlabel metal1 3751 -1896 3751 -1896 1 g2
rlabel metal1 4113 -171 4113 -171 1 y0d
rlabel metal1 4576 -1658 4576 -1658 1 y1d
rlabel metal1 5084 -1026 5084 -1026 1 e1
rlabel metal1 1607 358 1607 358 1 a1_f_1
rlabel metal1 756 208 756 208 1 vdd
rlabel metal1 1060 -51 1060 -51 1 gnd
rlabel metal1 3893 -225 3893 -225 1 lesser
rlabel metal1 5305 -1027 5305 -1027 1 equal
rlabel metal1 4087 -1762 4087 -1762 1 greater
<< end >>
