magic
tech scmos
timestamp 1699767830
<< nwell >>
rect -608 104 -570 120
rect -530 103 -492 119
rect -444 44 -406 60
rect -392 42 -351 60
rect -333 46 -295 62
rect -281 44 -240 62
rect -217 46 -179 62
rect -165 44 -124 62
rect -97 47 -59 63
rect -45 45 -4 63
rect 85 48 123 64
rect 137 46 178 64
rect 196 50 234 66
rect 248 48 289 66
rect 312 50 350 66
rect 364 48 405 66
rect 432 51 470 67
rect 484 49 525 67
rect -551 9 -513 25
rect -441 -158 -403 -142
rect -389 -160 -348 -142
rect -330 -156 -292 -140
rect -278 -158 -237 -140
rect -214 -156 -176 -140
rect -162 -158 -121 -140
rect -94 -155 -56 -139
rect -42 -157 -1 -139
rect 88 -154 126 -138
rect 140 -156 181 -138
rect 199 -152 237 -136
rect 251 -154 292 -136
rect 315 -152 353 -136
rect 367 -154 408 -136
rect 435 -151 473 -135
rect 487 -153 528 -135
rect -416 -335 -378 -319
rect -364 -337 -323 -319
rect -305 -333 -267 -317
rect -253 -335 -212 -317
rect -189 -333 -151 -317
rect -137 -335 -96 -317
rect -69 -332 -31 -316
rect -17 -334 24 -316
rect 113 -331 151 -315
rect 165 -333 206 -315
rect 224 -329 262 -313
rect 276 -331 317 -313
rect 340 -329 378 -313
rect 392 -331 433 -313
rect 460 -328 498 -312
rect 512 -330 553 -312
<< polysilicon >>
rect -596 114 -593 118
rect -585 114 -582 118
rect -518 113 -515 117
rect -507 113 -504 117
rect -596 103 -593 107
rect -596 83 -593 99
rect -585 95 -582 107
rect -518 102 -515 106
rect -585 83 -582 91
rect -518 82 -515 98
rect -507 94 -504 106
rect -507 82 -504 90
rect -596 71 -593 74
rect -585 71 -582 74
rect -518 70 -515 73
rect -507 70 -504 73
rect -432 54 -429 58
rect -421 54 -418 58
rect -374 54 -371 57
rect -321 56 -318 60
rect -310 56 -307 60
rect -263 56 -260 59
rect -205 56 -202 60
rect -194 56 -191 60
rect -147 56 -144 59
rect -85 57 -82 61
rect -74 57 -71 61
rect -27 57 -24 60
rect 97 58 100 62
rect 108 58 111 62
rect 155 58 158 61
rect 208 60 211 64
rect 219 60 222 64
rect 266 60 269 63
rect 324 60 327 64
rect 335 60 338 64
rect 382 60 385 63
rect 444 61 447 65
rect 455 61 458 65
rect 502 61 505 64
rect -432 43 -429 47
rect -432 23 -429 39
rect -421 35 -418 47
rect -374 34 -371 49
rect -321 45 -318 49
rect -421 23 -418 31
rect -539 19 -536 23
rect -528 19 -525 23
rect -374 15 -371 30
rect -321 25 -318 41
rect -310 37 -307 49
rect -263 36 -260 51
rect -205 45 -202 49
rect -310 25 -307 33
rect -263 17 -260 32
rect -205 25 -202 41
rect -194 37 -191 49
rect -147 36 -144 51
rect -85 46 -82 50
rect -194 25 -191 33
rect -539 8 -536 12
rect -539 -12 -536 4
rect -528 0 -525 12
rect -432 11 -429 14
rect -421 11 -418 14
rect -321 13 -318 16
rect -310 13 -307 16
rect -147 17 -144 32
rect -85 26 -82 42
rect -74 38 -71 50
rect -27 37 -24 52
rect 97 47 100 51
rect -74 26 -71 34
rect -27 18 -24 33
rect 97 27 100 43
rect 108 39 111 51
rect 155 38 158 53
rect 208 49 211 53
rect 108 27 111 35
rect 155 19 158 34
rect 208 29 211 45
rect 219 41 222 53
rect 266 40 269 55
rect 324 49 327 53
rect 219 29 222 37
rect 266 21 269 36
rect 324 29 327 45
rect 335 41 338 53
rect 382 40 385 55
rect 444 50 447 54
rect 335 29 338 37
rect -205 13 -202 16
rect -194 13 -191 16
rect -85 14 -82 17
rect -74 14 -71 17
rect 97 15 100 18
rect 108 15 111 18
rect 208 17 211 20
rect 219 17 222 20
rect 382 21 385 36
rect 444 30 447 46
rect 455 42 458 54
rect 502 41 505 56
rect 455 30 458 38
rect 502 22 505 37
rect 324 17 327 20
rect 335 17 338 20
rect 444 18 447 21
rect 455 18 458 21
rect -374 6 -371 10
rect -263 8 -260 12
rect -147 8 -144 12
rect -27 9 -24 13
rect 155 10 158 14
rect 266 12 269 16
rect 382 12 385 16
rect 502 13 505 17
rect -528 -12 -525 -4
rect -539 -24 -536 -21
rect -528 -24 -525 -21
rect -429 -148 -426 -144
rect -418 -148 -415 -144
rect -371 -148 -368 -145
rect -318 -146 -315 -142
rect -307 -146 -304 -142
rect -260 -146 -257 -143
rect -202 -146 -199 -142
rect -191 -146 -188 -142
rect -144 -146 -141 -143
rect -82 -145 -79 -141
rect -71 -145 -68 -141
rect -24 -145 -21 -142
rect 100 -144 103 -140
rect 111 -144 114 -140
rect 158 -144 161 -141
rect 211 -142 214 -138
rect 222 -142 225 -138
rect 269 -142 272 -139
rect 327 -142 330 -138
rect 338 -142 341 -138
rect 385 -142 388 -139
rect 447 -141 450 -137
rect 458 -141 461 -137
rect 505 -141 508 -138
rect -429 -159 -426 -155
rect -429 -179 -426 -163
rect -418 -167 -415 -155
rect -371 -168 -368 -153
rect -318 -157 -315 -153
rect -418 -179 -415 -171
rect -371 -187 -368 -172
rect -318 -177 -315 -161
rect -307 -165 -304 -153
rect -260 -166 -257 -151
rect -202 -157 -199 -153
rect -307 -177 -304 -169
rect -260 -185 -257 -170
rect -202 -177 -199 -161
rect -191 -165 -188 -153
rect -144 -166 -141 -151
rect -82 -156 -79 -152
rect -191 -177 -188 -169
rect -429 -191 -426 -188
rect -418 -191 -415 -188
rect -318 -189 -315 -186
rect -307 -189 -304 -186
rect -144 -185 -141 -170
rect -82 -176 -79 -160
rect -71 -164 -68 -152
rect -24 -165 -21 -150
rect 100 -155 103 -151
rect -71 -176 -68 -168
rect -24 -184 -21 -169
rect 100 -175 103 -159
rect 111 -163 114 -151
rect 158 -164 161 -149
rect 211 -153 214 -149
rect 111 -175 114 -167
rect 158 -183 161 -168
rect 211 -173 214 -157
rect 222 -161 225 -149
rect 269 -162 272 -147
rect 327 -153 330 -149
rect 222 -173 225 -165
rect 269 -181 272 -166
rect 327 -173 330 -157
rect 338 -161 341 -149
rect 385 -162 388 -147
rect 447 -152 450 -148
rect 338 -173 341 -165
rect -202 -189 -199 -186
rect -191 -189 -188 -186
rect -82 -188 -79 -185
rect -71 -188 -68 -185
rect 100 -187 103 -184
rect 111 -187 114 -184
rect 211 -185 214 -182
rect 222 -185 225 -182
rect 385 -181 388 -166
rect 447 -172 450 -156
rect 458 -160 461 -148
rect 505 -161 508 -146
rect 458 -172 461 -164
rect 505 -180 508 -165
rect 327 -185 330 -182
rect 338 -185 341 -182
rect 447 -184 450 -181
rect 458 -184 461 -181
rect -371 -196 -368 -192
rect -260 -194 -257 -190
rect -144 -194 -141 -190
rect -24 -193 -21 -189
rect 158 -192 161 -188
rect 269 -190 272 -186
rect 385 -190 388 -186
rect 505 -189 508 -185
rect -404 -325 -401 -321
rect -393 -325 -390 -321
rect -346 -325 -343 -322
rect -293 -323 -290 -319
rect -282 -323 -279 -319
rect -235 -323 -232 -320
rect -177 -323 -174 -319
rect -166 -323 -163 -319
rect -119 -323 -116 -320
rect -57 -322 -54 -318
rect -46 -322 -43 -318
rect 1 -322 4 -319
rect 125 -321 128 -317
rect 136 -321 139 -317
rect 183 -321 186 -318
rect 236 -319 239 -315
rect 247 -319 250 -315
rect 294 -319 297 -316
rect 352 -319 355 -315
rect 363 -319 366 -315
rect 410 -319 413 -316
rect 472 -318 475 -314
rect 483 -318 486 -314
rect 530 -318 533 -315
rect -404 -336 -401 -332
rect -404 -356 -401 -340
rect -393 -344 -390 -332
rect -346 -345 -343 -330
rect -293 -334 -290 -330
rect -393 -356 -390 -348
rect -346 -364 -343 -349
rect -293 -354 -290 -338
rect -282 -342 -279 -330
rect -235 -343 -232 -328
rect -177 -334 -174 -330
rect -282 -354 -279 -346
rect -235 -362 -232 -347
rect -177 -354 -174 -338
rect -166 -342 -163 -330
rect -119 -343 -116 -328
rect -57 -333 -54 -329
rect -166 -354 -163 -346
rect -404 -368 -401 -365
rect -393 -368 -390 -365
rect -293 -366 -290 -363
rect -282 -366 -279 -363
rect -119 -362 -116 -347
rect -57 -353 -54 -337
rect -46 -341 -43 -329
rect 1 -342 4 -327
rect 125 -332 128 -328
rect -46 -353 -43 -345
rect 1 -361 4 -346
rect 125 -352 128 -336
rect 136 -340 139 -328
rect 183 -341 186 -326
rect 236 -330 239 -326
rect 136 -352 139 -344
rect 183 -360 186 -345
rect 236 -350 239 -334
rect 247 -338 250 -326
rect 294 -339 297 -324
rect 352 -330 355 -326
rect 247 -350 250 -342
rect 294 -358 297 -343
rect 352 -350 355 -334
rect 363 -338 366 -326
rect 410 -339 413 -324
rect 472 -329 475 -325
rect 363 -350 366 -342
rect -177 -366 -174 -363
rect -166 -366 -163 -363
rect -57 -365 -54 -362
rect -46 -365 -43 -362
rect 125 -364 128 -361
rect 136 -364 139 -361
rect 236 -362 239 -359
rect 247 -362 250 -359
rect 410 -358 413 -343
rect 472 -349 475 -333
rect 483 -337 486 -325
rect 530 -338 533 -323
rect 483 -349 486 -341
rect 530 -357 533 -342
rect 352 -362 355 -359
rect 363 -362 366 -359
rect 472 -361 475 -358
rect 483 -361 486 -358
rect -346 -373 -343 -369
rect -235 -371 -232 -367
rect -119 -371 -116 -367
rect 1 -370 4 -366
rect 183 -369 186 -365
rect 294 -367 297 -363
rect 410 -367 413 -363
rect 530 -366 533 -362
<< ndiffusion >>
rect -598 79 -596 83
rect -602 74 -596 79
rect -593 74 -585 83
rect -582 79 -579 83
rect -575 79 -574 83
rect -582 74 -574 79
rect -520 78 -518 82
rect -524 73 -518 78
rect -515 73 -507 82
rect -504 78 -501 82
rect -497 78 -496 82
rect -504 73 -496 78
rect -434 19 -432 23
rect -438 14 -432 19
rect -429 14 -421 23
rect -418 19 -415 23
rect -411 19 -410 23
rect -418 14 -410 19
rect -323 21 -321 25
rect -327 16 -321 21
rect -318 16 -310 25
rect -307 21 -304 25
rect -300 21 -299 25
rect -307 16 -299 21
rect -207 21 -205 25
rect -377 10 -374 15
rect -371 10 -367 15
rect -266 12 -263 17
rect -260 12 -256 17
rect -211 16 -205 21
rect -202 16 -194 25
rect -191 21 -188 25
rect -184 21 -183 25
rect -191 16 -183 21
rect -87 22 -85 26
rect -91 17 -85 22
rect -82 17 -74 26
rect -71 22 -68 26
rect -64 22 -63 26
rect -71 17 -63 22
rect 95 23 97 27
rect 91 18 97 23
rect 100 18 108 27
rect 111 23 114 27
rect 118 23 119 27
rect 111 18 119 23
rect 206 25 208 29
rect 202 20 208 25
rect 211 20 219 29
rect 222 25 225 29
rect 229 25 230 29
rect 222 20 230 25
rect 322 25 324 29
rect -150 12 -147 17
rect -144 12 -140 17
rect -30 13 -27 18
rect -24 13 -20 18
rect 152 14 155 19
rect 158 14 162 19
rect 263 16 266 21
rect 269 16 273 21
rect 318 20 324 25
rect 327 20 335 29
rect 338 25 341 29
rect 345 25 346 29
rect 338 20 346 25
rect 442 26 444 30
rect 438 21 444 26
rect 447 21 455 30
rect 458 26 461 30
rect 465 26 466 30
rect 458 21 466 26
rect 379 16 382 21
rect 385 16 389 21
rect 499 17 502 22
rect 505 17 509 22
rect -541 -16 -539 -12
rect -545 -21 -539 -16
rect -536 -21 -528 -12
rect -525 -16 -522 -12
rect -518 -16 -517 -12
rect -525 -21 -517 -16
rect -431 -183 -429 -179
rect -435 -188 -429 -183
rect -426 -188 -418 -179
rect -415 -183 -412 -179
rect -408 -183 -407 -179
rect -415 -188 -407 -183
rect -320 -181 -318 -177
rect -324 -186 -318 -181
rect -315 -186 -307 -177
rect -304 -181 -301 -177
rect -297 -181 -296 -177
rect -304 -186 -296 -181
rect -204 -181 -202 -177
rect -374 -192 -371 -187
rect -368 -192 -364 -187
rect -263 -190 -260 -185
rect -257 -190 -253 -185
rect -208 -186 -202 -181
rect -199 -186 -191 -177
rect -188 -181 -185 -177
rect -181 -181 -180 -177
rect -188 -186 -180 -181
rect -84 -180 -82 -176
rect -88 -185 -82 -180
rect -79 -185 -71 -176
rect -68 -180 -65 -176
rect -61 -180 -60 -176
rect -68 -185 -60 -180
rect 98 -179 100 -175
rect 94 -184 100 -179
rect 103 -184 111 -175
rect 114 -179 117 -175
rect 121 -179 122 -175
rect 114 -184 122 -179
rect 209 -177 211 -173
rect 205 -182 211 -177
rect 214 -182 222 -173
rect 225 -177 228 -173
rect 232 -177 233 -173
rect 225 -182 233 -177
rect 325 -177 327 -173
rect -147 -190 -144 -185
rect -141 -190 -137 -185
rect -27 -189 -24 -184
rect -21 -189 -17 -184
rect 155 -188 158 -183
rect 161 -188 165 -183
rect 266 -186 269 -181
rect 272 -186 276 -181
rect 321 -182 327 -177
rect 330 -182 338 -173
rect 341 -177 344 -173
rect 348 -177 349 -173
rect 341 -182 349 -177
rect 445 -176 447 -172
rect 441 -181 447 -176
rect 450 -181 458 -172
rect 461 -176 464 -172
rect 468 -176 469 -172
rect 461 -181 469 -176
rect 382 -186 385 -181
rect 388 -186 392 -181
rect 502 -185 505 -180
rect 508 -185 512 -180
rect -406 -360 -404 -356
rect -410 -365 -404 -360
rect -401 -365 -393 -356
rect -390 -360 -387 -356
rect -383 -360 -382 -356
rect -390 -365 -382 -360
rect -295 -358 -293 -354
rect -299 -363 -293 -358
rect -290 -363 -282 -354
rect -279 -358 -276 -354
rect -272 -358 -271 -354
rect -279 -363 -271 -358
rect -179 -358 -177 -354
rect -349 -369 -346 -364
rect -343 -369 -339 -364
rect -238 -367 -235 -362
rect -232 -367 -228 -362
rect -183 -363 -177 -358
rect -174 -363 -166 -354
rect -163 -358 -160 -354
rect -156 -358 -155 -354
rect -163 -363 -155 -358
rect -59 -357 -57 -353
rect -63 -362 -57 -357
rect -54 -362 -46 -353
rect -43 -357 -40 -353
rect -36 -357 -35 -353
rect -43 -362 -35 -357
rect 123 -356 125 -352
rect 119 -361 125 -356
rect 128 -361 136 -352
rect 139 -356 142 -352
rect 146 -356 147 -352
rect 139 -361 147 -356
rect 234 -354 236 -350
rect 230 -359 236 -354
rect 239 -359 247 -350
rect 250 -354 253 -350
rect 257 -354 258 -350
rect 250 -359 258 -354
rect 350 -354 352 -350
rect -122 -367 -119 -362
rect -116 -367 -112 -362
rect -2 -366 1 -361
rect 4 -366 8 -361
rect 180 -365 183 -360
rect 186 -365 190 -360
rect 291 -363 294 -358
rect 297 -363 301 -358
rect 346 -359 352 -354
rect 355 -359 363 -350
rect 366 -354 369 -350
rect 373 -354 374 -350
rect 366 -359 374 -354
rect 470 -353 472 -349
rect 466 -358 472 -353
rect 475 -358 483 -349
rect 486 -353 489 -349
rect 493 -353 494 -349
rect 486 -358 494 -353
rect 407 -363 410 -358
rect 413 -363 417 -358
rect 527 -362 530 -357
rect 533 -362 537 -357
<< pdiffusion >>
rect -599 110 -596 114
rect -603 107 -596 110
rect -593 110 -590 114
rect -586 110 -585 114
rect -593 107 -585 110
rect -582 110 -579 114
rect -582 107 -575 110
rect -521 109 -518 113
rect -525 106 -518 109
rect -515 109 -512 113
rect -508 109 -507 113
rect -515 106 -507 109
rect -504 109 -501 113
rect -504 106 -497 109
rect -435 50 -432 54
rect -439 47 -432 50
rect -429 50 -426 54
rect -422 50 -421 54
rect -429 47 -421 50
rect -418 50 -415 54
rect -418 47 -411 50
rect -378 49 -374 54
rect -371 49 -367 54
rect -363 49 -361 54
rect -324 52 -321 56
rect -328 49 -321 52
rect -318 52 -315 56
rect -311 52 -310 56
rect -318 49 -310 52
rect -307 52 -304 56
rect -307 49 -300 52
rect -267 51 -263 56
rect -260 51 -256 56
rect -252 51 -250 56
rect -208 52 -205 56
rect -542 15 -539 19
rect -546 12 -539 15
rect -536 15 -533 19
rect -529 15 -528 19
rect -536 12 -528 15
rect -525 15 -522 19
rect -525 12 -518 15
rect -212 49 -205 52
rect -202 52 -199 56
rect -195 52 -194 56
rect -202 49 -194 52
rect -191 52 -188 56
rect -191 49 -184 52
rect -151 51 -147 56
rect -144 51 -140 56
rect -136 51 -134 56
rect -88 53 -85 57
rect -92 50 -85 53
rect -82 53 -79 57
rect -75 53 -74 57
rect -82 50 -74 53
rect -71 53 -68 57
rect -71 50 -64 53
rect -31 52 -27 57
rect -24 52 -20 57
rect -16 52 -14 57
rect 94 54 97 58
rect 90 51 97 54
rect 100 54 103 58
rect 107 54 108 58
rect 100 51 108 54
rect 111 54 114 58
rect 111 51 118 54
rect 151 53 155 58
rect 158 53 162 58
rect 166 53 168 58
rect 205 56 208 60
rect 201 53 208 56
rect 211 56 214 60
rect 218 56 219 60
rect 211 53 219 56
rect 222 56 225 60
rect 222 53 229 56
rect 262 55 266 60
rect 269 55 273 60
rect 277 55 279 60
rect 321 56 324 60
rect 317 53 324 56
rect 327 56 330 60
rect 334 56 335 60
rect 327 53 335 56
rect 338 56 341 60
rect 338 53 345 56
rect 378 55 382 60
rect 385 55 389 60
rect 393 55 395 60
rect 441 57 444 61
rect 437 54 444 57
rect 447 57 450 61
rect 454 57 455 61
rect 447 54 455 57
rect 458 57 461 61
rect 458 54 465 57
rect 498 56 502 61
rect 505 56 509 61
rect 513 56 515 61
rect -432 -152 -429 -148
rect -436 -155 -429 -152
rect -426 -152 -423 -148
rect -419 -152 -418 -148
rect -426 -155 -418 -152
rect -415 -152 -412 -148
rect -415 -155 -408 -152
rect -375 -153 -371 -148
rect -368 -153 -364 -148
rect -360 -153 -358 -148
rect -321 -150 -318 -146
rect -325 -153 -318 -150
rect -315 -150 -312 -146
rect -308 -150 -307 -146
rect -315 -153 -307 -150
rect -304 -150 -301 -146
rect -304 -153 -297 -150
rect -264 -151 -260 -146
rect -257 -151 -253 -146
rect -249 -151 -247 -146
rect -205 -150 -202 -146
rect -209 -153 -202 -150
rect -199 -150 -196 -146
rect -192 -150 -191 -146
rect -199 -153 -191 -150
rect -188 -150 -185 -146
rect -188 -153 -181 -150
rect -148 -151 -144 -146
rect -141 -151 -137 -146
rect -133 -151 -131 -146
rect -85 -149 -82 -145
rect -89 -152 -82 -149
rect -79 -149 -76 -145
rect -72 -149 -71 -145
rect -79 -152 -71 -149
rect -68 -149 -65 -145
rect -68 -152 -61 -149
rect -28 -150 -24 -145
rect -21 -150 -17 -145
rect -13 -150 -11 -145
rect 97 -148 100 -144
rect 93 -151 100 -148
rect 103 -148 106 -144
rect 110 -148 111 -144
rect 103 -151 111 -148
rect 114 -148 117 -144
rect 114 -151 121 -148
rect 154 -149 158 -144
rect 161 -149 165 -144
rect 169 -149 171 -144
rect 208 -146 211 -142
rect 204 -149 211 -146
rect 214 -146 217 -142
rect 221 -146 222 -142
rect 214 -149 222 -146
rect 225 -146 228 -142
rect 225 -149 232 -146
rect 265 -147 269 -142
rect 272 -147 276 -142
rect 280 -147 282 -142
rect 324 -146 327 -142
rect 320 -149 327 -146
rect 330 -146 333 -142
rect 337 -146 338 -142
rect 330 -149 338 -146
rect 341 -146 344 -142
rect 341 -149 348 -146
rect 381 -147 385 -142
rect 388 -147 392 -142
rect 396 -147 398 -142
rect 444 -145 447 -141
rect 440 -148 447 -145
rect 450 -145 453 -141
rect 457 -145 458 -141
rect 450 -148 458 -145
rect 461 -145 464 -141
rect 461 -148 468 -145
rect 501 -146 505 -141
rect 508 -146 512 -141
rect 516 -146 518 -141
rect -407 -329 -404 -325
rect -411 -332 -404 -329
rect -401 -329 -398 -325
rect -394 -329 -393 -325
rect -401 -332 -393 -329
rect -390 -329 -387 -325
rect -390 -332 -383 -329
rect -350 -330 -346 -325
rect -343 -330 -339 -325
rect -335 -330 -333 -325
rect -296 -327 -293 -323
rect -300 -330 -293 -327
rect -290 -327 -287 -323
rect -283 -327 -282 -323
rect -290 -330 -282 -327
rect -279 -327 -276 -323
rect -279 -330 -272 -327
rect -239 -328 -235 -323
rect -232 -328 -228 -323
rect -224 -328 -222 -323
rect -180 -327 -177 -323
rect -184 -330 -177 -327
rect -174 -327 -171 -323
rect -167 -327 -166 -323
rect -174 -330 -166 -327
rect -163 -327 -160 -323
rect -163 -330 -156 -327
rect -123 -328 -119 -323
rect -116 -328 -112 -323
rect -108 -328 -106 -323
rect -60 -326 -57 -322
rect -64 -329 -57 -326
rect -54 -326 -51 -322
rect -47 -326 -46 -322
rect -54 -329 -46 -326
rect -43 -326 -40 -322
rect -43 -329 -36 -326
rect -3 -327 1 -322
rect 4 -327 8 -322
rect 12 -327 14 -322
rect 122 -325 125 -321
rect 118 -328 125 -325
rect 128 -325 131 -321
rect 135 -325 136 -321
rect 128 -328 136 -325
rect 139 -325 142 -321
rect 139 -328 146 -325
rect 179 -326 183 -321
rect 186 -326 190 -321
rect 194 -326 196 -321
rect 233 -323 236 -319
rect 229 -326 236 -323
rect 239 -323 242 -319
rect 246 -323 247 -319
rect 239 -326 247 -323
rect 250 -323 253 -319
rect 250 -326 257 -323
rect 290 -324 294 -319
rect 297 -324 301 -319
rect 305 -324 307 -319
rect 349 -323 352 -319
rect 345 -326 352 -323
rect 355 -323 358 -319
rect 362 -323 363 -319
rect 355 -326 363 -323
rect 366 -323 369 -319
rect 366 -326 373 -323
rect 406 -324 410 -319
rect 413 -324 417 -319
rect 421 -324 423 -319
rect 469 -322 472 -318
rect 465 -325 472 -322
rect 475 -322 478 -318
rect 482 -322 483 -318
rect 475 -325 483 -322
rect 486 -322 489 -318
rect 486 -325 493 -322
rect 526 -323 530 -318
rect 533 -323 537 -318
rect 541 -323 543 -318
<< metal1 >>
rect -593 124 -588 125
rect -603 123 -510 124
rect -603 120 -497 123
rect -603 114 -599 120
rect -579 114 -575 120
rect -525 119 -497 120
rect -525 113 -521 119
rect -501 113 -497 119
rect -590 103 -586 110
rect -610 99 -597 103
rect -590 100 -575 103
rect -512 102 -508 109
rect -604 95 -601 99
rect -579 97 -575 100
rect -531 98 -519 102
rect -512 99 -497 102
rect -604 91 -586 95
rect -579 94 -574 97
rect -527 94 -523 98
rect -501 96 -497 99
rect -501 94 -496 96
rect -579 90 -567 94
rect -527 90 -508 94
rect -501 91 -489 94
rect -579 83 -575 90
rect -602 70 -598 79
rect -602 67 -573 70
rect -593 65 -586 67
rect -570 0 -567 90
rect -501 82 -497 91
rect -524 69 -520 78
rect -524 66 -495 69
rect -513 64 -507 66
rect -492 40 -489 91
rect 75 78 422 82
rect -454 77 422 78
rect -454 73 80 77
rect -454 57 -449 73
rect -564 37 -489 40
rect -477 53 -449 57
rect -564 8 -560 37
rect -536 29 -529 32
rect -546 25 -518 29
rect -546 19 -542 25
rect -522 19 -518 25
rect -533 8 -529 15
rect -564 4 -540 8
rect -533 5 -518 8
rect -522 2 -518 5
rect -477 2 -473 53
rect -454 43 -449 53
rect -439 60 -379 64
rect -375 60 -350 64
rect -439 54 -435 60
rect -415 54 -411 60
rect -382 54 -379 60
rect -426 43 -422 50
rect -454 39 -433 43
rect -426 40 -411 43
rect -442 31 -422 35
rect -415 34 -411 40
rect -415 30 -375 34
rect -415 23 -411 30
rect -438 10 -434 19
rect -366 15 -363 49
rect -344 45 -339 73
rect -328 62 -268 66
rect -264 62 -239 66
rect -328 56 -324 62
rect -304 56 -300 62
rect -271 56 -268 62
rect -315 45 -311 52
rect -344 41 -322 45
rect -315 42 -300 45
rect -304 39 -300 42
rect -331 33 -311 37
rect -304 36 -299 39
rect -304 32 -264 36
rect -304 25 -300 32
rect -327 12 -323 21
rect -255 17 -252 51
rect -226 45 -221 73
rect -212 62 -152 66
rect -148 62 -123 66
rect -212 56 -208 62
rect -188 56 -184 62
rect -155 56 -152 62
rect -199 45 -195 52
rect -226 41 -206 45
rect -199 42 -184 45
rect -188 39 -184 42
rect -215 33 -195 37
rect -188 36 -183 39
rect -188 32 -148 36
rect -188 25 -184 32
rect -211 12 -207 21
rect -139 17 -136 51
rect -112 46 -107 73
rect -92 63 -32 67
rect -28 63 -3 67
rect -92 57 -88 63
rect -68 57 -64 63
rect -35 57 -32 63
rect -79 46 -75 53
rect -112 42 -86 46
rect -79 43 -64 46
rect -68 40 -64 43
rect -95 34 -75 38
rect -68 37 -63 40
rect -68 33 -28 37
rect -68 26 -64 33
rect -91 13 -87 22
rect -19 18 -16 52
rect 74 47 80 73
rect 90 64 150 68
rect 154 64 179 68
rect 90 58 94 64
rect 114 58 118 64
rect 147 58 150 64
rect 103 47 107 54
rect 74 43 96 47
rect 103 44 118 47
rect 87 35 107 39
rect 114 38 118 44
rect 114 34 154 38
rect 114 27 118 34
rect 91 14 95 23
rect 163 19 166 53
rect 185 49 190 77
rect 201 66 261 70
rect 265 66 290 70
rect 201 60 205 66
rect 225 60 229 66
rect 258 60 261 66
rect 214 49 218 56
rect 185 45 207 49
rect 214 46 229 49
rect 225 43 229 46
rect 198 37 218 41
rect 225 40 230 43
rect 225 36 265 40
rect 225 29 229 36
rect 202 16 206 25
rect 274 21 277 55
rect 303 49 308 77
rect 317 66 377 70
rect 381 66 406 70
rect 317 60 321 66
rect 341 60 345 66
rect 374 60 377 66
rect 330 49 334 56
rect 303 45 323 49
rect 330 46 345 49
rect 341 43 345 46
rect 314 37 334 41
rect 341 40 346 43
rect 341 36 381 40
rect 341 29 345 36
rect 318 16 322 25
rect 390 21 393 55
rect 417 50 422 77
rect 437 67 497 71
rect 501 67 526 71
rect 437 61 441 67
rect 461 61 465 67
rect 494 61 497 67
rect 450 50 454 57
rect 417 46 443 50
rect 450 47 465 50
rect 461 44 465 47
rect 434 38 454 42
rect 461 41 466 44
rect 461 37 501 41
rect 461 30 465 37
rect 438 17 442 26
rect 510 22 513 56
rect -438 7 -392 10
rect -382 7 -378 10
rect -327 9 -281 12
rect -271 9 -267 12
rect -211 9 -165 12
rect -155 9 -151 12
rect -91 10 -45 13
rect -35 10 -31 13
rect 91 11 137 14
rect 147 11 151 14
rect 202 13 248 16
rect 258 13 262 16
rect 318 13 364 16
rect 374 13 378 16
rect 438 14 484 17
rect 494 14 498 17
rect -410 4 -378 7
rect -299 6 -267 9
rect -183 6 -151 9
rect -63 7 -31 10
rect 119 8 151 11
rect 230 10 262 13
rect 346 10 378 13
rect 466 11 498 14
rect -570 -4 -529 0
rect -522 -2 -473 2
rect -522 -12 -518 -2
rect -545 -25 -541 -16
rect -545 -28 -516 -25
rect -534 -30 -526 -28
rect 78 -123 425 -120
rect -106 -124 425 -123
rect -451 -125 425 -124
rect -451 -127 83 -125
rect -451 -129 -104 -127
rect -451 -159 -446 -129
rect -436 -142 -376 -138
rect -372 -142 -347 -138
rect -436 -148 -432 -142
rect -412 -148 -408 -142
rect -379 -148 -376 -142
rect -423 -159 -419 -152
rect -451 -163 -430 -159
rect -423 -162 -408 -159
rect -439 -171 -419 -167
rect -412 -168 -408 -162
rect -412 -172 -372 -168
rect -412 -179 -408 -172
rect -435 -192 -431 -183
rect -363 -187 -360 -153
rect -341 -157 -336 -129
rect -325 -140 -265 -136
rect -261 -140 -236 -136
rect -325 -146 -321 -140
rect -301 -146 -297 -140
rect -268 -146 -265 -140
rect -312 -157 -308 -150
rect -341 -161 -319 -157
rect -312 -160 -297 -157
rect -301 -163 -297 -160
rect -328 -169 -308 -165
rect -301 -166 -296 -163
rect -301 -170 -261 -166
rect -301 -177 -297 -170
rect -324 -190 -320 -181
rect -252 -185 -249 -151
rect -223 -157 -218 -129
rect -209 -140 -149 -136
rect -145 -140 -120 -136
rect -209 -146 -205 -140
rect -185 -146 -181 -140
rect -152 -146 -149 -140
rect -196 -157 -192 -150
rect -223 -161 -203 -157
rect -196 -160 -181 -157
rect -185 -163 -181 -160
rect -212 -169 -192 -165
rect -185 -166 -180 -163
rect -185 -170 -145 -166
rect -185 -177 -181 -170
rect -208 -190 -204 -181
rect -136 -185 -133 -151
rect -109 -156 -104 -129
rect -89 -139 -29 -135
rect -25 -139 0 -135
rect -89 -145 -85 -139
rect -65 -145 -61 -139
rect -32 -145 -29 -139
rect -76 -156 -72 -149
rect -109 -160 -83 -156
rect -76 -159 -61 -156
rect -65 -162 -61 -159
rect -92 -168 -72 -164
rect -65 -165 -60 -162
rect -65 -169 -25 -165
rect -65 -176 -61 -169
rect -88 -189 -84 -180
rect -16 -184 -13 -150
rect 78 -155 83 -127
rect 93 -138 153 -134
rect 157 -138 182 -134
rect 93 -144 97 -138
rect 117 -144 121 -138
rect 150 -144 153 -138
rect 106 -155 110 -148
rect 78 -159 99 -155
rect 106 -158 121 -155
rect 90 -167 110 -163
rect 117 -164 121 -158
rect 117 -168 157 -164
rect 117 -175 121 -168
rect 94 -188 98 -179
rect 166 -183 169 -149
rect 188 -153 193 -125
rect 204 -136 264 -132
rect 268 -136 293 -132
rect 204 -142 208 -136
rect 228 -142 232 -136
rect 261 -142 264 -136
rect 217 -153 221 -146
rect 188 -157 210 -153
rect 217 -156 232 -153
rect 228 -159 232 -156
rect 201 -165 221 -161
rect 228 -162 233 -159
rect 228 -166 268 -162
rect 228 -173 232 -166
rect 205 -186 209 -177
rect 277 -181 280 -147
rect 306 -153 311 -125
rect 320 -136 380 -132
rect 384 -136 409 -132
rect 320 -142 324 -136
rect 344 -142 348 -136
rect 377 -142 380 -136
rect 333 -153 337 -146
rect 306 -157 326 -153
rect 333 -156 348 -153
rect 344 -159 348 -156
rect 317 -165 337 -161
rect 344 -162 349 -159
rect 344 -166 384 -162
rect 344 -173 348 -166
rect 321 -186 325 -177
rect 393 -181 396 -147
rect 420 -152 425 -125
rect 440 -135 500 -131
rect 504 -135 529 -131
rect 440 -141 444 -135
rect 464 -141 468 -135
rect 497 -141 500 -135
rect 453 -152 457 -145
rect 420 -156 446 -152
rect 453 -155 468 -152
rect 464 -158 468 -155
rect 437 -164 457 -160
rect 464 -161 469 -158
rect 464 -165 504 -161
rect 464 -172 468 -165
rect 441 -185 445 -176
rect 513 -180 516 -146
rect -435 -195 -389 -192
rect -379 -195 -375 -192
rect -324 -193 -278 -190
rect -268 -193 -264 -190
rect -208 -193 -162 -190
rect -152 -193 -148 -190
rect -88 -192 -42 -189
rect -32 -192 -28 -189
rect 94 -191 140 -188
rect 150 -191 154 -188
rect 205 -189 251 -186
rect 261 -189 265 -186
rect 321 -189 367 -186
rect 377 -189 381 -186
rect 441 -188 487 -185
rect 497 -188 501 -185
rect -407 -198 -375 -195
rect -296 -196 -264 -193
rect -180 -196 -148 -193
rect -60 -195 -28 -192
rect 122 -194 154 -191
rect 233 -192 265 -189
rect 349 -192 381 -189
rect 469 -191 501 -188
rect 103 -301 450 -297
rect -426 -302 450 -301
rect -426 -304 108 -302
rect -426 -306 -79 -304
rect -426 -336 -421 -306
rect -411 -319 -351 -315
rect -347 -319 -322 -315
rect -411 -325 -407 -319
rect -387 -325 -383 -319
rect -354 -325 -351 -319
rect -398 -336 -394 -329
rect -426 -340 -405 -336
rect -398 -339 -383 -336
rect -414 -348 -394 -344
rect -387 -345 -383 -339
rect -387 -349 -347 -345
rect -387 -356 -383 -349
rect -410 -369 -406 -360
rect -338 -364 -335 -330
rect -316 -334 -311 -306
rect -300 -317 -240 -313
rect -236 -317 -211 -313
rect -300 -323 -296 -317
rect -276 -323 -272 -317
rect -243 -323 -240 -317
rect -287 -334 -283 -327
rect -316 -338 -294 -334
rect -287 -337 -272 -334
rect -276 -340 -272 -337
rect -303 -346 -283 -342
rect -276 -343 -271 -340
rect -276 -347 -236 -343
rect -276 -354 -272 -347
rect -299 -367 -295 -358
rect -227 -362 -224 -328
rect -198 -334 -193 -306
rect -184 -317 -124 -313
rect -120 -317 -95 -313
rect -184 -323 -180 -317
rect -160 -323 -156 -317
rect -127 -323 -124 -317
rect -171 -334 -167 -327
rect -198 -338 -178 -334
rect -171 -337 -156 -334
rect -160 -340 -156 -337
rect -187 -346 -167 -342
rect -160 -343 -155 -340
rect -160 -347 -120 -343
rect -160 -354 -156 -347
rect -183 -367 -179 -358
rect -111 -362 -108 -328
rect -84 -333 -79 -306
rect -64 -316 -4 -312
rect 0 -316 25 -312
rect -64 -322 -60 -316
rect -40 -322 -36 -316
rect -7 -322 -4 -316
rect -51 -333 -47 -326
rect -84 -337 -58 -333
rect -51 -336 -36 -333
rect -40 -339 -36 -336
rect -67 -345 -47 -341
rect -40 -342 -35 -339
rect -40 -346 0 -342
rect -40 -353 -36 -346
rect -63 -366 -59 -357
rect 9 -361 12 -327
rect 103 -332 108 -304
rect 118 -315 178 -311
rect 182 -315 207 -311
rect 118 -321 122 -315
rect 142 -321 146 -315
rect 175 -321 178 -315
rect 131 -332 135 -325
rect 103 -336 124 -332
rect 131 -335 146 -332
rect 115 -344 135 -340
rect 142 -341 146 -335
rect 142 -345 182 -341
rect 142 -352 146 -345
rect 119 -365 123 -356
rect 191 -360 194 -326
rect 213 -330 218 -302
rect 229 -313 289 -309
rect 293 -313 318 -309
rect 229 -319 233 -313
rect 253 -319 257 -313
rect 286 -319 289 -313
rect 242 -330 246 -323
rect 213 -334 235 -330
rect 242 -333 257 -330
rect 253 -336 257 -333
rect 226 -342 246 -338
rect 253 -339 258 -336
rect 253 -343 293 -339
rect 253 -350 257 -343
rect 230 -363 234 -354
rect 302 -358 305 -324
rect 331 -330 336 -302
rect 345 -313 405 -309
rect 409 -313 434 -309
rect 345 -319 349 -313
rect 369 -319 373 -313
rect 402 -319 405 -313
rect 358 -330 362 -323
rect 331 -334 351 -330
rect 358 -333 373 -330
rect 369 -336 373 -333
rect 342 -342 362 -338
rect 369 -339 374 -336
rect 369 -343 409 -339
rect 369 -350 373 -343
rect 346 -363 350 -354
rect 418 -358 421 -324
rect 445 -329 450 -302
rect 465 -312 525 -308
rect 529 -312 554 -308
rect 465 -318 469 -312
rect 489 -318 493 -312
rect 522 -318 525 -312
rect 478 -329 482 -322
rect 445 -333 471 -329
rect 478 -332 493 -329
rect 489 -335 493 -332
rect 462 -341 482 -337
rect 489 -338 494 -335
rect 489 -342 529 -338
rect 489 -349 493 -342
rect 466 -362 470 -353
rect 538 -357 541 -323
rect -410 -372 -364 -369
rect -354 -372 -350 -369
rect -299 -370 -253 -367
rect -243 -370 -239 -367
rect -183 -370 -137 -367
rect -127 -370 -123 -367
rect -63 -369 -17 -366
rect -7 -369 -3 -366
rect 119 -368 165 -365
rect 175 -368 179 -365
rect 230 -366 276 -363
rect 286 -366 290 -363
rect 346 -366 392 -363
rect 402 -366 406 -363
rect 466 -365 512 -362
rect 522 -365 526 -362
rect -382 -375 -350 -372
rect -271 -373 -239 -370
rect -155 -373 -123 -370
rect -35 -372 -3 -369
rect 147 -371 179 -368
rect 258 -369 290 -366
rect 374 -369 406 -366
rect 494 -368 526 -365
<< ntransistor >>
rect -596 74 -593 83
rect -585 74 -582 83
rect -518 73 -515 82
rect -507 73 -504 82
rect -432 14 -429 23
rect -421 14 -418 23
rect -321 16 -318 25
rect -310 16 -307 25
rect -374 10 -371 15
rect -263 12 -260 17
rect -205 16 -202 25
rect -194 16 -191 25
rect -85 17 -82 26
rect -74 17 -71 26
rect 97 18 100 27
rect 108 18 111 27
rect 208 20 211 29
rect 219 20 222 29
rect -147 12 -144 17
rect -27 13 -24 18
rect 155 14 158 19
rect 266 16 269 21
rect 324 20 327 29
rect 335 20 338 29
rect 444 21 447 30
rect 455 21 458 30
rect 382 16 385 21
rect 502 17 505 22
rect -539 -21 -536 -12
rect -528 -21 -525 -12
rect -429 -188 -426 -179
rect -418 -188 -415 -179
rect -318 -186 -315 -177
rect -307 -186 -304 -177
rect -371 -192 -368 -187
rect -260 -190 -257 -185
rect -202 -186 -199 -177
rect -191 -186 -188 -177
rect -82 -185 -79 -176
rect -71 -185 -68 -176
rect 100 -184 103 -175
rect 111 -184 114 -175
rect 211 -182 214 -173
rect 222 -182 225 -173
rect -144 -190 -141 -185
rect -24 -189 -21 -184
rect 158 -188 161 -183
rect 269 -186 272 -181
rect 327 -182 330 -173
rect 338 -182 341 -173
rect 447 -181 450 -172
rect 458 -181 461 -172
rect 385 -186 388 -181
rect 505 -185 508 -180
rect -404 -365 -401 -356
rect -393 -365 -390 -356
rect -293 -363 -290 -354
rect -282 -363 -279 -354
rect -346 -369 -343 -364
rect -235 -367 -232 -362
rect -177 -363 -174 -354
rect -166 -363 -163 -354
rect -57 -362 -54 -353
rect -46 -362 -43 -353
rect 125 -361 128 -352
rect 136 -361 139 -352
rect 236 -359 239 -350
rect 247 -359 250 -350
rect -119 -367 -116 -362
rect 1 -366 4 -361
rect 183 -365 186 -360
rect 294 -363 297 -358
rect 352 -359 355 -350
rect 363 -359 366 -350
rect 472 -358 475 -349
rect 483 -358 486 -349
rect 410 -363 413 -358
rect 530 -362 533 -357
<< ptransistor >>
rect -596 107 -593 114
rect -585 107 -582 114
rect -518 106 -515 113
rect -507 106 -504 113
rect -432 47 -429 54
rect -421 47 -418 54
rect -374 49 -371 54
rect -321 49 -318 56
rect -310 49 -307 56
rect -263 51 -260 56
rect -539 12 -536 19
rect -528 12 -525 19
rect -205 49 -202 56
rect -194 49 -191 56
rect -147 51 -144 56
rect -85 50 -82 57
rect -74 50 -71 57
rect -27 52 -24 57
rect 97 51 100 58
rect 108 51 111 58
rect 155 53 158 58
rect 208 53 211 60
rect 219 53 222 60
rect 266 55 269 60
rect 324 53 327 60
rect 335 53 338 60
rect 382 55 385 60
rect 444 54 447 61
rect 455 54 458 61
rect 502 56 505 61
rect -429 -155 -426 -148
rect -418 -155 -415 -148
rect -371 -153 -368 -148
rect -318 -153 -315 -146
rect -307 -153 -304 -146
rect -260 -151 -257 -146
rect -202 -153 -199 -146
rect -191 -153 -188 -146
rect -144 -151 -141 -146
rect -82 -152 -79 -145
rect -71 -152 -68 -145
rect -24 -150 -21 -145
rect 100 -151 103 -144
rect 111 -151 114 -144
rect 158 -149 161 -144
rect 211 -149 214 -142
rect 222 -149 225 -142
rect 269 -147 272 -142
rect 327 -149 330 -142
rect 338 -149 341 -142
rect 385 -147 388 -142
rect 447 -148 450 -141
rect 458 -148 461 -141
rect 505 -146 508 -141
rect -404 -332 -401 -325
rect -393 -332 -390 -325
rect -346 -330 -343 -325
rect -293 -330 -290 -323
rect -282 -330 -279 -323
rect -235 -328 -232 -323
rect -177 -330 -174 -323
rect -166 -330 -163 -323
rect -119 -328 -116 -323
rect -57 -329 -54 -322
rect -46 -329 -43 -322
rect 1 -327 4 -322
rect 125 -328 128 -321
rect 136 -328 139 -321
rect 183 -326 186 -321
rect 236 -326 239 -319
rect 247 -326 250 -319
rect 294 -324 297 -319
rect 352 -326 355 -319
rect 363 -326 366 -319
rect 410 -324 413 -319
rect 472 -325 475 -318
rect 483 -325 486 -318
rect 530 -323 533 -318
<< polycontact >>
rect -597 99 -593 103
rect -519 98 -515 102
rect -586 91 -582 95
rect -508 90 -504 94
rect -433 39 -429 43
rect -422 31 -418 35
rect -322 41 -318 45
rect -375 30 -371 34
rect -311 33 -307 37
rect -206 41 -202 45
rect -264 32 -260 36
rect -195 33 -191 37
rect -86 42 -82 46
rect -148 32 -144 36
rect -540 4 -536 8
rect -75 34 -71 38
rect 96 43 100 47
rect -28 33 -24 37
rect 107 35 111 39
rect 207 45 211 49
rect 154 34 158 38
rect 218 37 222 41
rect 323 45 327 49
rect 265 36 269 40
rect 334 37 338 41
rect 443 46 447 50
rect 381 36 385 40
rect 454 38 458 42
rect 501 37 505 41
rect -529 -4 -525 0
rect -430 -163 -426 -159
rect -419 -171 -415 -167
rect -319 -161 -315 -157
rect -372 -172 -368 -168
rect -308 -169 -304 -165
rect -203 -161 -199 -157
rect -261 -170 -257 -166
rect -192 -169 -188 -165
rect -83 -160 -79 -156
rect -145 -170 -141 -166
rect -72 -168 -68 -164
rect 99 -159 103 -155
rect -25 -169 -21 -165
rect 110 -167 114 -163
rect 210 -157 214 -153
rect 157 -168 161 -164
rect 221 -165 225 -161
rect 326 -157 330 -153
rect 268 -166 272 -162
rect 337 -165 341 -161
rect 446 -156 450 -152
rect 384 -166 388 -162
rect 457 -164 461 -160
rect 504 -165 508 -161
rect -405 -340 -401 -336
rect -394 -348 -390 -344
rect -294 -338 -290 -334
rect -347 -349 -343 -345
rect -283 -346 -279 -342
rect -178 -338 -174 -334
rect -236 -347 -232 -343
rect -167 -346 -163 -342
rect -58 -337 -54 -333
rect -120 -347 -116 -343
rect -47 -345 -43 -341
rect 124 -336 128 -332
rect 0 -346 4 -342
rect 135 -344 139 -340
rect 235 -334 239 -330
rect 182 -345 186 -341
rect 246 -342 250 -338
rect 351 -334 355 -330
rect 293 -343 297 -339
rect 362 -342 366 -338
rect 471 -333 475 -329
rect 409 -343 413 -339
rect 482 -341 486 -337
rect 529 -342 533 -338
<< ndcontact >>
rect -602 79 -598 83
rect -579 79 -575 83
rect -524 78 -520 82
rect -501 78 -497 82
rect -438 19 -434 23
rect -415 19 -411 23
rect -327 21 -323 25
rect -304 21 -300 25
rect -211 21 -207 25
rect -382 10 -377 15
rect -367 10 -363 15
rect -271 12 -266 17
rect -256 12 -252 17
rect -188 21 -184 25
rect -91 22 -87 26
rect -68 22 -64 26
rect 91 23 95 27
rect 114 23 118 27
rect 202 25 206 29
rect 225 25 229 29
rect 318 25 322 29
rect -155 12 -150 17
rect -140 12 -136 17
rect -35 13 -30 18
rect -20 13 -16 18
rect 147 14 152 19
rect 162 14 166 19
rect 258 16 263 21
rect 273 16 277 21
rect 341 25 345 29
rect 438 26 442 30
rect 461 26 465 30
rect 374 16 379 21
rect 389 16 393 21
rect 494 17 499 22
rect 509 17 513 22
rect -545 -16 -541 -12
rect -522 -16 -518 -12
rect -435 -183 -431 -179
rect -412 -183 -408 -179
rect -324 -181 -320 -177
rect -301 -181 -297 -177
rect -208 -181 -204 -177
rect -379 -192 -374 -187
rect -364 -192 -360 -187
rect -268 -190 -263 -185
rect -253 -190 -249 -185
rect -185 -181 -181 -177
rect -88 -180 -84 -176
rect -65 -180 -61 -176
rect 94 -179 98 -175
rect 117 -179 121 -175
rect 205 -177 209 -173
rect 228 -177 232 -173
rect 321 -177 325 -173
rect -152 -190 -147 -185
rect -137 -190 -133 -185
rect -32 -189 -27 -184
rect -17 -189 -13 -184
rect 150 -188 155 -183
rect 165 -188 169 -183
rect 261 -186 266 -181
rect 276 -186 280 -181
rect 344 -177 348 -173
rect 441 -176 445 -172
rect 464 -176 468 -172
rect 377 -186 382 -181
rect 392 -186 396 -181
rect 497 -185 502 -180
rect 512 -185 516 -180
rect -410 -360 -406 -356
rect -387 -360 -383 -356
rect -299 -358 -295 -354
rect -276 -358 -272 -354
rect -183 -358 -179 -354
rect -354 -369 -349 -364
rect -339 -369 -335 -364
rect -243 -367 -238 -362
rect -228 -367 -224 -362
rect -160 -358 -156 -354
rect -63 -357 -59 -353
rect -40 -357 -36 -353
rect 119 -356 123 -352
rect 142 -356 146 -352
rect 230 -354 234 -350
rect 253 -354 257 -350
rect 346 -354 350 -350
rect -127 -367 -122 -362
rect -112 -367 -108 -362
rect -7 -366 -2 -361
rect 8 -366 12 -361
rect 175 -365 180 -360
rect 190 -365 194 -360
rect 286 -363 291 -358
rect 301 -363 305 -358
rect 369 -354 373 -350
rect 466 -353 470 -349
rect 489 -353 493 -349
rect 402 -363 407 -358
rect 417 -363 421 -358
rect 522 -362 527 -357
rect 537 -362 541 -357
<< pdcontact >>
rect -603 110 -599 114
rect -590 110 -586 114
rect -579 110 -575 114
rect -525 109 -521 113
rect -512 109 -508 113
rect -501 109 -497 113
rect -439 50 -435 54
rect -426 50 -422 54
rect -415 50 -411 54
rect -382 49 -378 54
rect -367 49 -363 54
rect -328 52 -324 56
rect -315 52 -311 56
rect -304 52 -300 56
rect -271 51 -267 56
rect -256 51 -252 56
rect -212 52 -208 56
rect -546 15 -542 19
rect -533 15 -529 19
rect -522 15 -518 19
rect -199 52 -195 56
rect -188 52 -184 56
rect -155 51 -151 56
rect -140 51 -136 56
rect -92 53 -88 57
rect -79 53 -75 57
rect -68 53 -64 57
rect -35 52 -31 57
rect -20 52 -16 57
rect 90 54 94 58
rect 103 54 107 58
rect 114 54 118 58
rect 147 53 151 58
rect 162 53 166 58
rect 201 56 205 60
rect 214 56 218 60
rect 225 56 229 60
rect 258 55 262 60
rect 273 55 277 60
rect 317 56 321 60
rect 330 56 334 60
rect 341 56 345 60
rect 374 55 378 60
rect 389 55 393 60
rect 437 57 441 61
rect 450 57 454 61
rect 461 57 465 61
rect 494 56 498 61
rect 509 56 513 61
rect -436 -152 -432 -148
rect -423 -152 -419 -148
rect -412 -152 -408 -148
rect -379 -153 -375 -148
rect -364 -153 -360 -148
rect -325 -150 -321 -146
rect -312 -150 -308 -146
rect -301 -150 -297 -146
rect -268 -151 -264 -146
rect -253 -151 -249 -146
rect -209 -150 -205 -146
rect -196 -150 -192 -146
rect -185 -150 -181 -146
rect -152 -151 -148 -146
rect -137 -151 -133 -146
rect -89 -149 -85 -145
rect -76 -149 -72 -145
rect -65 -149 -61 -145
rect -32 -150 -28 -145
rect -17 -150 -13 -145
rect 93 -148 97 -144
rect 106 -148 110 -144
rect 117 -148 121 -144
rect 150 -149 154 -144
rect 165 -149 169 -144
rect 204 -146 208 -142
rect 217 -146 221 -142
rect 228 -146 232 -142
rect 261 -147 265 -142
rect 276 -147 280 -142
rect 320 -146 324 -142
rect 333 -146 337 -142
rect 344 -146 348 -142
rect 377 -147 381 -142
rect 392 -147 396 -142
rect 440 -145 444 -141
rect 453 -145 457 -141
rect 464 -145 468 -141
rect 497 -146 501 -141
rect 512 -146 516 -141
rect -411 -329 -407 -325
rect -398 -329 -394 -325
rect -387 -329 -383 -325
rect -354 -330 -350 -325
rect -339 -330 -335 -325
rect -300 -327 -296 -323
rect -287 -327 -283 -323
rect -276 -327 -272 -323
rect -243 -328 -239 -323
rect -228 -328 -224 -323
rect -184 -327 -180 -323
rect -171 -327 -167 -323
rect -160 -327 -156 -323
rect -127 -328 -123 -323
rect -112 -328 -108 -323
rect -64 -326 -60 -322
rect -51 -326 -47 -322
rect -40 -326 -36 -322
rect -7 -327 -3 -322
rect 8 -327 12 -322
rect 118 -325 122 -321
rect 131 -325 135 -321
rect 142 -325 146 -321
rect 175 -326 179 -321
rect 190 -326 194 -321
rect 229 -323 233 -319
rect 242 -323 246 -319
rect 253 -323 257 -319
rect 286 -324 290 -319
rect 301 -324 305 -319
rect 345 -323 349 -319
rect 358 -323 362 -319
rect 369 -323 373 -319
rect 402 -324 406 -319
rect 417 -324 421 -319
rect 465 -322 469 -318
rect 478 -322 482 -318
rect 489 -322 493 -318
rect 522 -323 526 -318
rect 537 -323 541 -318
<< nsubstratencontact >>
rect -379 60 -375 64
rect -268 62 -264 66
rect -152 62 -148 66
rect -32 63 -28 67
rect 150 64 154 68
rect 261 66 265 70
rect 377 66 381 70
rect 497 67 501 71
rect -376 -142 -372 -138
rect -265 -140 -261 -136
rect -149 -140 -145 -136
rect -29 -139 -25 -135
rect 153 -138 157 -134
rect 264 -136 268 -132
rect 380 -136 384 -132
rect 500 -135 504 -131
rect -351 -319 -347 -315
rect -240 -317 -236 -313
rect -124 -317 -120 -313
rect -4 -316 0 -312
rect 178 -315 182 -311
rect 289 -313 293 -309
rect 405 -313 409 -309
rect 525 -312 529 -308
<< labels >>
rlabel metal1 130 11 130 11 1 gnd
rlabel metal1 241 13 241 13 1 gnd
rlabel metal1 357 13 357 13 1 gnd
rlabel metal1 477 14 477 14 1 gnd
rlabel metal1 90 37 90 37 1 B0
rlabel metal1 165 35 165 35 1 b1_f_0
rlabel metal1 201 38 201 38 1 B1
rlabel metal1 276 38 276 38 1 b1_f_1
rlabel metal1 317 38 317 38 1 B2
rlabel metal1 391 37 391 37 1 b1_f_2
rlabel metal1 438 40 438 40 1 B3
rlabel metal1 511 38 511 38 1 b1_f_3
rlabel metal1 478 69 478 69 1 vdd
rlabel metal1 130 67 130 67 1 vdd
rlabel metal1 242 68 242 68 1 vdd
rlabel metal1 358 69 358 69 1 vdd
rlabel metal1 -396 -195 -396 -195 1 gnd
rlabel metal1 -285 -193 -285 -193 1 gnd
rlabel metal1 -169 -193 -169 -193 1 gnd
rlabel metal1 -49 -192 -49 -192 1 gnd
rlabel metal1 -437 -169 -437 -169 1 A0
rlabel metal1 -324 -167 -324 -167 1 A1
rlabel metal1 -208 -168 -208 -168 1 A2
rlabel metal1 -89 -165 -89 -165 1 A3
rlabel metal1 -399 -140 -399 -140 1 vdd
rlabel metal1 -287 -138 -287 -138 1 vdd
rlabel metal1 -175 -137 -175 -137 1 vdd
rlabel metal1 -50 -137 -50 -137 1 vdd
rlabel metal1 -371 -372 -371 -372 1 gnd
rlabel metal1 -260 -370 -260 -370 1 gnd
rlabel metal1 -144 -370 -144 -370 1 gnd
rlabel metal1 -24 -369 -24 -369 1 gnd
rlabel metal1 -412 -346 -412 -346 1 A0
rlabel metal1 -299 -344 -299 -344 1 A1
rlabel metal1 -183 -345 -183 -345 1 A2
rlabel metal1 -64 -342 -64 -342 1 A3
rlabel metal1 -374 -317 -374 -317 1 vdd
rlabel metal1 -262 -315 -262 -315 1 vdd
rlabel metal1 -150 -314 -150 -314 1 vdd
rlabel metal1 -25 -314 -25 -314 1 vdd
rlabel metal1 -425 -324 -425 -324 1 D3
rlabel metal1 -450 -138 -449 -138 3 D2
rlabel metal1 -549 121 -549 122 5 vdd
rlabel metal1 -533 29 -533 29 1 vdd
rlabel metal1 -591 68 -591 68 1 gnd
rlabel metal1 -509 66 -509 66 1 gnd
rlabel metal1 -530 -28 -530 -28 1 gnd
rlabel metal1 -609 101 -609 101 3 D0
rlabel metal1 -530 100 -530 100 1 D1
rlabel metal1 -53 65 -53 65 1 vdd
rlabel metal1 -178 65 -178 65 1 vdd
rlabel metal1 -290 64 -290 64 1 vdd
rlabel metal1 -402 62 -402 62 1 vdd
rlabel metal1 -17 33 -17 33 1 a1_f_3
rlabel metal1 -137 34 -137 34 1 a1_f_2
rlabel metal1 -254 33 -254 33 1 a1_f_1
rlabel metal1 -365 32 -365 32 1 a1_f_0
rlabel metal1 -92 37 -92 37 1 A3
rlabel metal1 -211 34 -211 34 1 A2
rlabel metal1 -327 35 -327 35 1 A1
rlabel metal1 -440 33 -440 33 1 A0
rlabel metal1 -52 10 -52 10 1 gnd
rlabel metal1 -172 9 -172 9 1 gnd
rlabel metal1 -288 9 -288 9 1 gnd
rlabel metal1 -399 7 -399 7 1 gnd
rlabel metal1 -361 -170 -361 -170 1 a2_f_0
rlabel metal1 -250 -168 -250 -168 1 a2_f_1
rlabel metal1 -135 -168 -135 -168 1 a2_f_2
rlabel metal1 -15 -169 -15 -169 1 a2_f_3
rlabel metal1 -336 -346 -336 -346 1 a3_f_0
rlabel metal1 -226 -344 -226 -344 1 a3_f_1
rlabel metal1 -109 -344 -109 -344 1 a3_f_2
rlabel metal1 10 -344 10 -344 1 a3_f_3
rlabel metal1 386 -310 386 -310 1 vdd
rlabel metal1 270 -311 270 -311 1 vdd
rlabel metal1 158 -312 158 -312 1 vdd
rlabel metal1 506 -310 506 -310 1 vdd
rlabel metal1 466 -339 466 -339 1 B3
rlabel metal1 345 -341 345 -341 1 B2
rlabel metal1 229 -341 229 -341 1 B1
rlabel metal1 118 -342 118 -342 1 B0
rlabel metal1 505 -365 505 -365 1 gnd
rlabel metal1 385 -366 385 -366 1 gnd
rlabel metal1 269 -366 269 -366 1 gnd
rlabel metal1 158 -368 158 -368 1 gnd
rlabel metal1 361 -133 361 -133 1 vdd
rlabel metal1 245 -134 245 -134 1 vdd
rlabel metal1 133 -135 133 -135 1 vdd
rlabel metal1 481 -133 481 -133 1 vdd
rlabel metal1 441 -162 441 -162 1 B3
rlabel metal1 320 -164 320 -164 1 B2
rlabel metal1 204 -164 204 -164 1 B1
rlabel metal1 93 -165 93 -165 1 B0
rlabel metal1 480 -188 480 -188 1 gnd
rlabel metal1 360 -189 360 -189 1 gnd
rlabel metal1 244 -189 244 -189 1 gnd
rlabel metal1 133 -191 133 -191 1 gnd
rlabel metal1 -452 70 -452 70 1 deff
rlabel metal1 167 -166 167 -166 1 b2_f_0
rlabel metal1 278 -163 278 -163 1 b2_f_1
rlabel metal1 394 -163 394 -163 1 b2_f_2
rlabel metal1 514 -163 514 -163 1 b2_f_3
rlabel metal1 192 -344 192 -344 1 b3_f_0
rlabel metal1 303 -341 303 -341 1 b3_f_1
rlabel metal1 419 -340 419 -340 1 b3_f_2
rlabel metal1 539 -341 539 -341 1 b3_f_3
<< end >>
