.subckt NAND node_a node_b node_out vdd gnd

    Mn1 node_out node_a node_y gnd CMOSN W = {wn1} L = {ln1}
    + AS = {5*wn1*LAMBDA} PS = {10*LAMBDA + 2*wn1} AD = {5*wn1*LAMBDA} PD = {10*LAMBDA + 2*wn1}

    Mn2 node_y node_b gnd gnd CMOSN W = {wn2} L = {ln2}
    + AS = {5*wn2*LAMBDA} PS = {10*LAMBDA + 2*wn2} AD = {5*wn2*LAMBDA} PD = {10*LAMBDA + 2*wn2}

    Mp1 node_out node_a vdd vdd CMOSP W = {wp1} L = {lp1}
    + AS = {5*wp1*LAMBDA} PS = {10*LAMBDA + 2*wp1} AD = {5*wp1*LAMBDA} PD = {10*LAMBDA + 2*wp1}

    Mp2 node_out node_b vdd vdd CMOSP W = {wp2} L = {lp2}
    + AS = {5*wp2*LAMBDA} PS = {10*LAMBDA + 2*wp2} AD = {5*wp2*LAMBDA} PD = {10*LAMBDA + 2*wp2}

.ends NAND


   * AS: Short-channel drain current coefficient for strong inversion (AS)
   * PS: Short-channel source current coefficient for strong inversion (PS)
   * AD: Short-channel drain current coefficient for moderate inversion (AD)
   * PD: Short-channel source current coefficient for moderate inversion (PD)	
   
