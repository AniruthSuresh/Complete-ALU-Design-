
.subckt And4bit a3 a2 a1 a0 b3 b2 b1 b0 y3 y2 y1 y0 node_x gnd

	X1 a0 b0 y0 node_x gnd AND
	X2 a1 b1 y1 node_x gnd AND
	X3 a2 b2 y2 node_x gnd AND
	X4 a3 b3 y3 node_x gnd AND

.ends And4bit




