magic
tech scmos
timestamp 1699617909
<< nwell >>
rect -7 14 31 30
<< polysilicon >>
rect 5 24 8 28
rect 16 24 19 28
rect 5 13 8 17
rect 5 -7 8 9
rect 16 5 19 17
rect 16 -7 19 1
rect 5 -19 8 -16
rect 16 -19 19 -16
<< ndiffusion >>
rect 3 -11 5 -7
rect -1 -16 5 -11
rect 8 -16 16 -7
rect 19 -11 22 -7
rect 26 -11 27 -7
rect 19 -16 27 -11
<< pdiffusion >>
rect 2 20 5 24
rect -2 17 5 20
rect 8 20 11 24
rect 15 20 16 24
rect 8 17 16 20
rect 19 20 22 24
rect 19 17 26 20
<< metal1 >>
rect 8 34 13 35
rect -2 30 26 34
rect -2 24 2 30
rect 22 24 26 30
rect 11 13 15 20
rect -1 9 4 13
rect 11 10 26 13
rect 22 7 26 10
rect -1 1 15 5
rect 22 3 27 7
rect 22 -7 26 3
rect -1 -20 3 -11
rect -1 -23 28 -20
<< ntransistor >>
rect 5 -16 8 -7
rect 16 -16 19 -7
<< ptransistor >>
rect 5 17 8 24
rect 16 17 19 24
<< polycontact >>
rect 4 9 8 13
rect 15 1 19 5
<< ndcontact >>
rect -1 -11 3 -7
rect 22 -11 26 -7
<< pdcontact >>
rect -2 20 2 24
rect 11 20 15 24
rect 22 20 26 24
<< labels >>
rlabel metal1 -1 11 -1 11 1 A
rlabel metal1 -1 3 -1 3 1 B
rlabel metal1 27 5 27 5 7 out
rlabel metal1 10 35 10 35 5 vdd
rlabel metal1 28 -21 28 -21 8 gnd
<< end >>
