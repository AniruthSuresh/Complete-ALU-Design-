

.subckt XNOR node_a node_b node_out node_x gnd

	X1 node_a node_b node_d node_x gnd NAND
	X2 node_a node_d node_c node_x gnd NAND
	X3 node_d node_b node_e node_x gnd NAND
	X4 node_c node_e node_f node_x gnd NAND
	X5 node_f node_f node_out node_x gnd NAND
	
	*X1 node_a node_b node_c node_x gnd XOR
	*X2 node_c node_out node_x gnd NOT


.ends XNOR



