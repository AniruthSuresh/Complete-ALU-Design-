magic
tech scmos
timestamp 1699793617
<< nwell >>
rect 667 661 705 677
rect 745 660 783 676
rect 724 566 762 582
rect 885 534 923 550
rect 963 533 1001 549
rect 1173 495 1214 513
rect 942 439 980 455
rect 680 385 718 401
rect 758 384 796 400
rect 737 290 775 306
rect -94 51 -53 69
rect 71 51 112 69
rect 248 52 289 70
rect 423 51 464 69
rect 821 6 862 24
rect 911 -9 991 14
rect 1069 5 1110 23
rect 1312 14 1353 32
rect 1159 -10 1239 13
rect 1402 -1 1482 22
rect 1581 19 1622 37
rect 1671 4 1751 27
rect -43 -66 -5 -50
rect 9 -68 50 -50
rect 128 -61 166 -45
rect 180 -63 221 -45
rect 321 -65 359 -49
rect 373 -67 414 -49
rect 502 -61 540 -45
rect 554 -63 595 -45
rect 1160 -122 1198 -106
rect 1212 -124 1253 -106
rect 1380 -142 1418 -126
rect 1432 -144 1473 -126
rect 1536 -134 1574 -118
rect 1588 -136 1629 -118
rect 89 -205 127 -189
rect 141 -207 182 -189
rect 939 -237 977 -221
rect 991 -239 1032 -221
rect 2090 -359 2128 -343
rect 2142 -361 2183 -343
rect 2307 -359 2345 -343
rect 2359 -361 2400 -343
rect 93 -403 131 -387
rect 145 -405 186 -387
rect 1280 -406 1318 -390
rect 952 -423 990 -407
rect 1004 -425 1045 -407
rect 1332 -408 1373 -390
rect -69 -580 -28 -562
rect 96 -580 137 -562
rect 273 -579 314 -561
rect 448 -580 489 -562
rect -18 -697 20 -681
rect 34 -699 75 -681
rect 153 -692 191 -676
rect 205 -694 246 -676
rect 346 -696 384 -680
rect 398 -698 439 -680
rect 527 -692 565 -676
rect 579 -694 620 -676
rect 739 -893 777 -877
rect 817 -894 855 -878
rect 796 -988 834 -972
rect 1084 -1003 1122 -987
rect 1162 -1004 1200 -988
rect 1635 -992 1676 -974
rect 1141 -1098 1179 -1082
rect 749 -1137 787 -1121
rect 827 -1138 865 -1122
rect 806 -1232 844 -1216
<< polysilicon >>
rect 679 671 682 675
rect 690 671 693 675
rect 757 670 760 674
rect 768 670 771 674
rect 679 660 682 664
rect 679 640 682 656
rect 690 652 693 664
rect 757 659 760 663
rect 690 640 693 648
rect 757 639 760 655
rect 768 651 771 663
rect 768 639 771 647
rect 679 628 682 631
rect 690 628 693 631
rect 757 627 760 630
rect 768 627 771 630
rect 736 576 739 580
rect 747 576 750 580
rect 736 565 739 569
rect 736 545 739 561
rect 747 557 750 569
rect 747 545 750 553
rect 897 544 900 548
rect 908 544 911 548
rect 975 543 978 547
rect 986 543 989 547
rect 736 533 739 536
rect 747 533 750 536
rect 897 533 900 537
rect 897 513 900 529
rect 908 525 911 537
rect 975 532 978 536
rect 908 513 911 521
rect 975 512 978 528
rect 986 524 989 536
rect 986 512 989 520
rect 897 501 900 504
rect 908 501 911 504
rect 1191 507 1194 510
rect 975 500 978 503
rect 986 500 989 503
rect 1191 487 1194 502
rect 1191 468 1194 483
rect 1191 459 1194 463
rect 954 449 957 453
rect 965 449 968 453
rect 954 438 957 442
rect 954 418 957 434
rect 965 430 968 442
rect 965 418 968 426
rect 954 406 957 409
rect 965 406 968 409
rect 692 395 695 399
rect 703 395 706 399
rect 770 394 773 398
rect 781 394 784 398
rect 692 384 695 388
rect 692 364 695 380
rect 703 376 706 388
rect 770 383 773 387
rect 703 364 706 372
rect 770 363 773 379
rect 781 375 784 387
rect 781 363 784 371
rect 692 352 695 355
rect 703 352 706 355
rect 770 351 773 354
rect 781 351 784 354
rect 749 300 752 304
rect 760 300 763 304
rect 749 289 752 293
rect 749 269 752 285
rect 760 281 763 293
rect 760 269 763 277
rect 749 257 752 260
rect 760 257 763 260
rect -76 63 -73 66
rect 89 63 92 66
rect 266 64 269 67
rect 441 63 444 66
rect -76 43 -73 58
rect 89 43 92 58
rect 266 44 269 59
rect 441 43 444 58
rect 1663 47 1699 49
rect -76 24 -73 39
rect 89 24 92 39
rect 266 25 269 40
rect 441 24 444 39
rect 1394 42 1430 44
rect 903 34 939 36
rect -76 15 -73 19
rect 89 15 92 19
rect 266 16 269 20
rect 441 15 444 19
rect 839 18 842 21
rect 839 -2 842 13
rect 839 -21 842 -6
rect 839 -30 842 -26
rect 903 -43 905 34
rect 918 5 920 7
rect 937 5 939 34
rect 1151 33 1187 35
rect 1087 17 1090 20
rect 962 5 964 7
rect 981 5 983 7
rect 918 -12 920 0
rect 937 -2 939 0
rect 962 -12 964 0
rect 918 -14 939 -12
rect 918 -26 920 -23
rect 937 -26 939 -14
rect 963 -16 964 -12
rect 962 -26 964 -16
rect 981 -26 983 0
rect 1087 -3 1090 12
rect 992 -15 998 -13
rect 918 -43 920 -31
rect 937 -39 939 -31
rect 962 -33 964 -31
rect 981 -39 983 -31
rect 937 -41 983 -39
rect 996 -43 998 -15
rect 1087 -22 1090 -7
rect 1087 -31 1090 -27
rect 903 -45 998 -43
rect 1151 -44 1153 33
rect 1166 4 1168 6
rect 1185 4 1187 33
rect 1330 26 1333 29
rect 1330 6 1333 21
rect 1210 4 1212 6
rect 1229 4 1231 6
rect 1166 -13 1168 -1
rect 1185 -3 1187 -1
rect 1210 -13 1212 -1
rect 1166 -15 1187 -13
rect 1166 -27 1168 -24
rect 1185 -27 1187 -15
rect 1211 -17 1212 -13
rect 1210 -27 1212 -17
rect 1229 -27 1231 -1
rect 1330 -13 1333 2
rect 1240 -16 1246 -14
rect 1166 -44 1168 -32
rect 1185 -40 1187 -32
rect 1210 -34 1212 -32
rect 1229 -40 1231 -32
rect 1185 -42 1231 -40
rect 1244 -44 1246 -16
rect 1330 -22 1333 -18
rect 1394 -35 1396 42
rect 1409 13 1411 15
rect 1428 13 1430 42
rect 1599 31 1602 34
rect 1453 13 1455 15
rect 1472 13 1474 15
rect 1599 11 1602 26
rect 1409 -4 1411 8
rect 1428 6 1430 8
rect 1453 -4 1455 8
rect 1409 -6 1430 -4
rect 1409 -18 1411 -15
rect 1428 -18 1430 -6
rect 1454 -8 1455 -4
rect 1453 -18 1455 -8
rect 1472 -18 1474 8
rect 1483 -7 1489 -5
rect 1409 -35 1411 -23
rect 1428 -31 1430 -23
rect 1453 -25 1455 -23
rect 1472 -31 1474 -23
rect 1428 -33 1474 -31
rect 1487 -35 1489 -7
rect 1599 -8 1602 7
rect 1599 -17 1602 -13
rect 1663 -30 1665 47
rect 1678 18 1680 20
rect 1697 18 1699 47
rect 1722 18 1724 20
rect 1741 18 1743 20
rect 1678 1 1680 13
rect 1697 11 1699 13
rect 1722 1 1724 13
rect 1678 -1 1699 1
rect 1678 -13 1680 -10
rect 1697 -13 1699 -1
rect 1723 -3 1724 1
rect 1722 -13 1724 -3
rect 1741 -13 1743 13
rect 1752 -2 1758 0
rect 1678 -30 1680 -18
rect 1697 -26 1699 -18
rect 1722 -20 1724 -18
rect 1741 -26 1743 -18
rect 1697 -28 1743 -26
rect 1756 -30 1758 -2
rect 1663 -32 1758 -30
rect 1394 -37 1489 -35
rect 140 -51 143 -47
rect 151 -51 154 -47
rect 198 -51 201 -48
rect 1151 -46 1246 -44
rect 514 -51 517 -47
rect 525 -51 528 -47
rect 572 -51 575 -48
rect -31 -56 -28 -52
rect -20 -56 -17 -52
rect 27 -56 30 -53
rect 333 -55 336 -51
rect 344 -55 347 -51
rect 391 -55 394 -52
rect -31 -67 -28 -63
rect -31 -87 -28 -71
rect -20 -75 -17 -63
rect 27 -76 30 -61
rect 140 -62 143 -58
rect -20 -87 -17 -79
rect 27 -95 30 -80
rect 140 -82 143 -66
rect 151 -70 154 -58
rect 198 -71 201 -56
rect 333 -66 336 -62
rect 151 -82 154 -74
rect 198 -90 201 -75
rect 333 -86 336 -70
rect 344 -74 347 -62
rect 391 -75 394 -60
rect 514 -62 517 -58
rect 344 -86 347 -78
rect 140 -94 143 -91
rect 151 -94 154 -91
rect 391 -94 394 -79
rect 514 -82 517 -66
rect 525 -70 528 -58
rect 572 -71 575 -56
rect 525 -82 528 -74
rect 572 -90 575 -75
rect 514 -94 517 -91
rect 525 -94 528 -91
rect -31 -99 -28 -96
rect -20 -99 -17 -96
rect 198 -99 201 -95
rect 333 -98 336 -95
rect 344 -98 347 -95
rect 572 -99 575 -95
rect 27 -104 30 -100
rect 391 -103 394 -99
rect 1172 -112 1175 -108
rect 1183 -112 1186 -108
rect 1230 -112 1233 -109
rect 1172 -123 1175 -119
rect 1172 -143 1175 -127
rect 1183 -131 1186 -119
rect 1230 -132 1233 -117
rect 1548 -124 1551 -120
rect 1559 -124 1562 -120
rect 1606 -124 1609 -121
rect 1392 -132 1395 -128
rect 1403 -132 1406 -128
rect 1450 -132 1453 -129
rect 1183 -143 1186 -135
rect 1230 -151 1233 -136
rect 1548 -135 1551 -131
rect 1392 -143 1395 -139
rect 1172 -155 1175 -152
rect 1183 -155 1186 -152
rect 1230 -160 1233 -156
rect 1392 -163 1395 -147
rect 1403 -151 1406 -139
rect 1450 -152 1453 -137
rect 1403 -163 1406 -155
rect 1548 -155 1551 -139
rect 1559 -143 1562 -131
rect 1606 -144 1609 -129
rect 1559 -155 1562 -147
rect 1450 -171 1453 -156
rect 1606 -163 1609 -148
rect 1548 -167 1551 -164
rect 1559 -167 1562 -164
rect 1392 -175 1395 -172
rect 1403 -175 1406 -172
rect 1606 -172 1609 -168
rect 1450 -180 1453 -176
rect 101 -195 104 -191
rect 112 -195 115 -191
rect 159 -195 162 -192
rect 101 -206 104 -202
rect 101 -226 104 -210
rect 112 -214 115 -202
rect 159 -215 162 -200
rect 112 -226 115 -218
rect 159 -234 162 -219
rect 951 -227 954 -223
rect 962 -227 965 -223
rect 1009 -227 1012 -224
rect 101 -238 104 -235
rect 112 -238 115 -235
rect 951 -238 954 -234
rect 159 -243 162 -239
rect 951 -258 954 -242
rect 962 -246 965 -234
rect 1009 -247 1012 -232
rect 962 -258 965 -250
rect 1009 -266 1012 -251
rect 951 -270 954 -267
rect 962 -270 965 -267
rect 1009 -275 1012 -271
rect 2102 -349 2105 -345
rect 2113 -349 2116 -345
rect 2160 -349 2163 -346
rect 2319 -349 2322 -345
rect 2330 -349 2333 -345
rect 2377 -349 2380 -346
rect 2102 -360 2105 -356
rect 2102 -380 2105 -364
rect 2113 -368 2116 -356
rect 2160 -369 2163 -354
rect 2319 -360 2322 -356
rect 2113 -380 2116 -372
rect 105 -393 108 -389
rect 116 -393 119 -389
rect 2160 -388 2163 -373
rect 2319 -380 2322 -364
rect 2330 -368 2333 -356
rect 2377 -369 2380 -354
rect 2330 -380 2333 -372
rect 163 -393 166 -390
rect 2102 -392 2105 -389
rect 2113 -392 2116 -389
rect 1292 -396 1295 -392
rect 1303 -396 1306 -392
rect 2377 -388 2380 -373
rect 2319 -392 2322 -389
rect 2330 -392 2333 -389
rect 1350 -396 1353 -393
rect 105 -404 108 -400
rect 105 -424 108 -408
rect 116 -412 119 -400
rect 163 -413 166 -398
rect 2160 -397 2163 -393
rect 2377 -397 2380 -393
rect 1292 -407 1295 -403
rect 964 -413 967 -409
rect 975 -413 978 -409
rect 1022 -413 1025 -410
rect 116 -424 119 -416
rect 163 -432 166 -417
rect 964 -424 967 -420
rect 105 -436 108 -433
rect 116 -436 119 -433
rect 163 -441 166 -437
rect 964 -444 967 -428
rect 975 -432 978 -420
rect 1022 -433 1025 -418
rect 1292 -427 1295 -411
rect 1303 -415 1306 -403
rect 1350 -416 1353 -401
rect 1303 -427 1306 -419
rect 975 -444 978 -436
rect 1350 -435 1353 -420
rect 1022 -452 1025 -437
rect 1292 -439 1295 -436
rect 1303 -439 1306 -436
rect 1350 -444 1353 -440
rect 964 -456 967 -453
rect 975 -456 978 -453
rect 1022 -461 1025 -457
rect -51 -568 -48 -565
rect 114 -568 117 -565
rect 291 -567 294 -564
rect 466 -568 469 -565
rect -51 -588 -48 -573
rect 114 -588 117 -573
rect 291 -587 294 -572
rect 466 -588 469 -573
rect -51 -607 -48 -592
rect 114 -607 117 -592
rect 291 -606 294 -591
rect 466 -607 469 -592
rect -51 -616 -48 -612
rect 114 -616 117 -612
rect 291 -615 294 -611
rect 466 -616 469 -612
rect 165 -682 168 -678
rect 176 -682 179 -678
rect 223 -682 226 -679
rect 539 -682 542 -678
rect 550 -682 553 -678
rect 597 -682 600 -679
rect -6 -687 -3 -683
rect 5 -687 8 -683
rect 52 -687 55 -684
rect 358 -686 361 -682
rect 369 -686 372 -682
rect 416 -686 419 -683
rect -6 -698 -3 -694
rect -6 -718 -3 -702
rect 5 -706 8 -694
rect 52 -707 55 -692
rect 165 -693 168 -689
rect 5 -718 8 -710
rect 52 -726 55 -711
rect 165 -713 168 -697
rect 176 -701 179 -689
rect 223 -702 226 -687
rect 358 -697 361 -693
rect 176 -713 179 -705
rect 223 -721 226 -706
rect 358 -717 361 -701
rect 369 -705 372 -693
rect 416 -706 419 -691
rect 539 -693 542 -689
rect 369 -717 372 -709
rect 165 -725 168 -722
rect 176 -725 179 -722
rect 416 -725 419 -710
rect 539 -713 542 -697
rect 550 -701 553 -689
rect 597 -702 600 -687
rect 550 -713 553 -705
rect 597 -721 600 -706
rect 539 -725 542 -722
rect 550 -725 553 -722
rect -6 -730 -3 -727
rect 5 -730 8 -727
rect 223 -730 226 -726
rect 358 -729 361 -726
rect 369 -729 372 -726
rect 597 -730 600 -726
rect 52 -735 55 -731
rect 416 -734 419 -730
rect 751 -883 754 -879
rect 762 -883 765 -879
rect 829 -884 832 -880
rect 840 -884 843 -880
rect 751 -894 754 -890
rect 751 -914 754 -898
rect 762 -902 765 -890
rect 829 -895 832 -891
rect 762 -914 765 -906
rect 829 -915 832 -899
rect 840 -903 843 -891
rect 840 -915 843 -907
rect 751 -926 754 -923
rect 762 -926 765 -923
rect 829 -927 832 -924
rect 840 -927 843 -924
rect 808 -978 811 -974
rect 819 -978 822 -974
rect 1653 -980 1656 -977
rect 808 -989 811 -985
rect 808 -1009 811 -993
rect 819 -997 822 -985
rect 1096 -993 1099 -989
rect 1107 -993 1110 -989
rect 1174 -994 1177 -990
rect 1185 -994 1188 -990
rect 819 -1009 822 -1001
rect 1096 -1004 1099 -1000
rect 808 -1021 811 -1018
rect 819 -1021 822 -1018
rect 1096 -1024 1099 -1008
rect 1107 -1012 1110 -1000
rect 1653 -1000 1656 -985
rect 1174 -1005 1177 -1001
rect 1107 -1024 1110 -1016
rect 1174 -1025 1177 -1009
rect 1185 -1013 1188 -1001
rect 1185 -1025 1188 -1017
rect 1653 -1019 1656 -1004
rect 1096 -1036 1099 -1033
rect 1107 -1036 1110 -1033
rect 1653 -1028 1656 -1024
rect 1174 -1037 1177 -1034
rect 1185 -1037 1188 -1034
rect 1153 -1088 1156 -1084
rect 1164 -1088 1167 -1084
rect 1153 -1099 1156 -1095
rect 1153 -1119 1156 -1103
rect 1164 -1107 1167 -1095
rect 1164 -1119 1167 -1111
rect 761 -1127 764 -1123
rect 772 -1127 775 -1123
rect 839 -1128 842 -1124
rect 850 -1128 853 -1124
rect 761 -1138 764 -1134
rect 761 -1158 764 -1142
rect 772 -1146 775 -1134
rect 1153 -1131 1156 -1128
rect 1164 -1131 1167 -1128
rect 839 -1139 842 -1135
rect 772 -1158 775 -1150
rect 839 -1159 842 -1143
rect 850 -1147 853 -1135
rect 850 -1159 853 -1151
rect 761 -1170 764 -1167
rect 772 -1170 775 -1167
rect 839 -1171 842 -1168
rect 850 -1171 853 -1168
rect 818 -1222 821 -1218
rect 829 -1222 832 -1218
rect 818 -1233 821 -1229
rect 818 -1253 821 -1237
rect 829 -1241 832 -1229
rect 829 -1253 832 -1245
rect 818 -1265 821 -1262
rect 829 -1265 832 -1262
<< ndiffusion >>
rect 677 636 679 640
rect 673 631 679 636
rect 682 631 690 640
rect 693 636 696 640
rect 700 636 701 640
rect 693 631 701 636
rect 755 635 757 639
rect 751 630 757 635
rect 760 630 768 639
rect 771 635 774 639
rect 778 635 779 639
rect 771 630 779 635
rect 734 541 736 545
rect 730 536 736 541
rect 739 536 747 545
rect 750 541 753 545
rect 757 541 758 545
rect 750 536 758 541
rect 895 509 897 513
rect 891 504 897 509
rect 900 504 908 513
rect 911 509 914 513
rect 918 509 919 513
rect 911 504 919 509
rect 973 508 975 512
rect 969 503 975 508
rect 978 503 986 512
rect 989 508 992 512
rect 996 508 997 512
rect 989 503 997 508
rect 1188 463 1191 468
rect 1194 463 1198 468
rect 952 414 954 418
rect 948 409 954 414
rect 957 409 965 418
rect 968 414 971 418
rect 975 414 976 418
rect 968 409 976 414
rect 690 360 692 364
rect 686 355 692 360
rect 695 355 703 364
rect 706 360 709 364
rect 713 360 714 364
rect 706 355 714 360
rect 768 359 770 363
rect 764 354 770 359
rect 773 354 781 363
rect 784 359 787 363
rect 791 359 792 363
rect 784 354 792 359
rect 747 265 749 269
rect 743 260 749 265
rect 752 260 760 269
rect 763 265 766 269
rect 770 265 771 269
rect 763 260 771 265
rect -79 19 -76 24
rect -73 19 -69 24
rect 86 19 89 24
rect 92 19 96 24
rect 263 20 266 25
rect 269 20 273 25
rect 438 19 441 24
rect 444 19 448 24
rect 836 -26 839 -21
rect 842 -26 846 -21
rect 915 -27 918 -26
rect 917 -31 918 -27
rect 920 -27 924 -26
rect 934 -27 937 -26
rect 920 -31 922 -27
rect 936 -31 937 -27
rect 939 -27 945 -26
rect 939 -31 941 -27
rect 957 -27 962 -26
rect 961 -31 962 -27
rect 964 -27 967 -26
rect 976 -27 981 -26
rect 964 -31 966 -27
rect 980 -31 981 -27
rect 983 -27 987 -26
rect 983 -31 985 -27
rect 1084 -27 1087 -22
rect 1090 -27 1094 -22
rect 1163 -28 1166 -27
rect 1165 -32 1166 -28
rect 1168 -28 1172 -27
rect 1182 -28 1185 -27
rect 1168 -32 1170 -28
rect 1184 -32 1185 -28
rect 1187 -28 1193 -27
rect 1187 -32 1189 -28
rect 1205 -28 1210 -27
rect 1209 -32 1210 -28
rect 1212 -28 1215 -27
rect 1224 -28 1229 -27
rect 1212 -32 1214 -28
rect 1228 -32 1229 -28
rect 1231 -28 1235 -27
rect 1231 -32 1233 -28
rect 1327 -18 1330 -13
rect 1333 -18 1337 -13
rect 1406 -19 1409 -18
rect 1408 -23 1409 -19
rect 1411 -19 1415 -18
rect 1425 -19 1428 -18
rect 1411 -23 1413 -19
rect 1427 -23 1428 -19
rect 1430 -19 1436 -18
rect 1430 -23 1432 -19
rect 1448 -19 1453 -18
rect 1452 -23 1453 -19
rect 1455 -19 1458 -18
rect 1467 -19 1472 -18
rect 1455 -23 1457 -19
rect 1471 -23 1472 -19
rect 1474 -19 1478 -18
rect 1474 -23 1476 -19
rect 1596 -13 1599 -8
rect 1602 -13 1606 -8
rect 1675 -14 1678 -13
rect 1677 -18 1678 -14
rect 1680 -14 1684 -13
rect 1694 -14 1697 -13
rect 1680 -18 1682 -14
rect 1696 -18 1697 -14
rect 1699 -14 1705 -13
rect 1699 -18 1701 -14
rect 1717 -14 1722 -13
rect 1721 -18 1722 -14
rect 1724 -14 1727 -13
rect 1736 -14 1741 -13
rect 1724 -18 1726 -14
rect 1740 -18 1741 -14
rect 1743 -14 1747 -13
rect 1743 -18 1745 -14
rect -33 -91 -31 -87
rect -37 -96 -31 -91
rect -28 -96 -20 -87
rect -17 -91 -14 -87
rect -10 -91 -9 -87
rect -17 -96 -9 -91
rect 138 -86 140 -82
rect 134 -91 140 -86
rect 143 -91 151 -82
rect 154 -86 157 -82
rect 161 -86 162 -82
rect 154 -91 162 -86
rect 331 -90 333 -86
rect 195 -95 198 -90
rect 201 -95 205 -90
rect 327 -95 333 -90
rect 336 -95 344 -86
rect 347 -90 350 -86
rect 354 -90 355 -86
rect 347 -95 355 -90
rect 512 -86 514 -82
rect 508 -91 514 -86
rect 517 -91 525 -82
rect 528 -86 531 -82
rect 535 -86 536 -82
rect 528 -91 536 -86
rect 24 -100 27 -95
rect 30 -100 34 -95
rect 388 -99 391 -94
rect 394 -99 398 -94
rect 569 -95 572 -90
rect 575 -95 579 -90
rect 1170 -147 1172 -143
rect 1166 -152 1172 -147
rect 1175 -152 1183 -143
rect 1186 -147 1189 -143
rect 1193 -147 1194 -143
rect 1186 -152 1194 -147
rect 1227 -156 1230 -151
rect 1233 -156 1237 -151
rect 1390 -167 1392 -163
rect 1386 -172 1392 -167
rect 1395 -172 1403 -163
rect 1406 -167 1409 -163
rect 1413 -167 1414 -163
rect 1406 -172 1414 -167
rect 1546 -159 1548 -155
rect 1542 -164 1548 -159
rect 1551 -164 1559 -155
rect 1562 -159 1565 -155
rect 1569 -159 1570 -155
rect 1562 -164 1570 -159
rect 1603 -168 1606 -163
rect 1609 -168 1613 -163
rect 1447 -176 1450 -171
rect 1453 -176 1457 -171
rect 99 -230 101 -226
rect 95 -235 101 -230
rect 104 -235 112 -226
rect 115 -230 118 -226
rect 122 -230 123 -226
rect 115 -235 123 -230
rect 156 -239 159 -234
rect 162 -239 166 -234
rect 949 -262 951 -258
rect 945 -267 951 -262
rect 954 -267 962 -258
rect 965 -262 968 -258
rect 972 -262 973 -258
rect 965 -267 973 -262
rect 1006 -271 1009 -266
rect 1012 -271 1016 -266
rect 2100 -384 2102 -380
rect 2096 -389 2102 -384
rect 2105 -389 2113 -380
rect 2116 -384 2119 -380
rect 2123 -384 2124 -380
rect 2116 -389 2124 -384
rect 2317 -384 2319 -380
rect 2157 -393 2160 -388
rect 2163 -393 2167 -388
rect 2313 -389 2319 -384
rect 2322 -389 2330 -380
rect 2333 -384 2336 -380
rect 2340 -384 2341 -380
rect 2333 -389 2341 -384
rect 2374 -393 2377 -388
rect 2380 -393 2384 -388
rect 103 -428 105 -424
rect 99 -433 105 -428
rect 108 -433 116 -424
rect 119 -428 122 -424
rect 126 -428 127 -424
rect 119 -433 127 -428
rect 160 -437 163 -432
rect 166 -437 170 -432
rect 1290 -431 1292 -427
rect 1286 -436 1292 -431
rect 1295 -436 1303 -427
rect 1306 -431 1309 -427
rect 1313 -431 1314 -427
rect 1306 -436 1314 -431
rect 962 -448 964 -444
rect 958 -453 964 -448
rect 967 -453 975 -444
rect 978 -448 981 -444
rect 985 -448 986 -444
rect 978 -453 986 -448
rect 1347 -440 1350 -435
rect 1353 -440 1357 -435
rect 1019 -457 1022 -452
rect 1025 -457 1029 -452
rect -54 -612 -51 -607
rect -48 -612 -44 -607
rect 111 -612 114 -607
rect 117 -612 121 -607
rect 288 -611 291 -606
rect 294 -611 298 -606
rect 463 -612 466 -607
rect 469 -612 473 -607
rect -8 -722 -6 -718
rect -12 -727 -6 -722
rect -3 -727 5 -718
rect 8 -722 11 -718
rect 15 -722 16 -718
rect 8 -727 16 -722
rect 163 -717 165 -713
rect 159 -722 165 -717
rect 168 -722 176 -713
rect 179 -717 182 -713
rect 186 -717 187 -713
rect 179 -722 187 -717
rect 356 -721 358 -717
rect 220 -726 223 -721
rect 226 -726 230 -721
rect 352 -726 358 -721
rect 361 -726 369 -717
rect 372 -721 375 -717
rect 379 -721 380 -717
rect 372 -726 380 -721
rect 537 -717 539 -713
rect 533 -722 539 -717
rect 542 -722 550 -713
rect 553 -717 556 -713
rect 560 -717 561 -713
rect 553 -722 561 -717
rect 49 -731 52 -726
rect 55 -731 59 -726
rect 413 -730 416 -725
rect 419 -730 423 -725
rect 594 -726 597 -721
rect 600 -726 604 -721
rect 749 -918 751 -914
rect 745 -923 751 -918
rect 754 -923 762 -914
rect 765 -918 768 -914
rect 772 -918 773 -914
rect 765 -923 773 -918
rect 827 -919 829 -915
rect 823 -924 829 -919
rect 832 -924 840 -915
rect 843 -919 846 -915
rect 850 -919 851 -915
rect 843 -924 851 -919
rect 806 -1013 808 -1009
rect 802 -1018 808 -1013
rect 811 -1018 819 -1009
rect 822 -1013 825 -1009
rect 829 -1013 830 -1009
rect 822 -1018 830 -1013
rect 1094 -1028 1096 -1024
rect 1090 -1033 1096 -1028
rect 1099 -1033 1107 -1024
rect 1110 -1028 1113 -1024
rect 1117 -1028 1118 -1024
rect 1650 -1024 1653 -1019
rect 1656 -1024 1660 -1019
rect 1110 -1033 1118 -1028
rect 1172 -1029 1174 -1025
rect 1168 -1034 1174 -1029
rect 1177 -1034 1185 -1025
rect 1188 -1029 1191 -1025
rect 1195 -1029 1196 -1025
rect 1188 -1034 1196 -1029
rect 1151 -1123 1153 -1119
rect 1147 -1128 1153 -1123
rect 1156 -1128 1164 -1119
rect 1167 -1123 1170 -1119
rect 1174 -1123 1175 -1119
rect 1167 -1128 1175 -1123
rect 759 -1162 761 -1158
rect 755 -1167 761 -1162
rect 764 -1167 772 -1158
rect 775 -1162 778 -1158
rect 782 -1162 783 -1158
rect 775 -1167 783 -1162
rect 837 -1163 839 -1159
rect 833 -1168 839 -1163
rect 842 -1168 850 -1159
rect 853 -1163 856 -1159
rect 860 -1163 861 -1159
rect 853 -1168 861 -1163
rect 816 -1257 818 -1253
rect 812 -1262 818 -1257
rect 821 -1262 829 -1253
rect 832 -1257 835 -1253
rect 839 -1257 840 -1253
rect 832 -1262 840 -1257
<< pdiffusion >>
rect 676 667 679 671
rect 672 664 679 667
rect 682 667 685 671
rect 689 667 690 671
rect 682 664 690 667
rect 693 667 696 671
rect 693 664 700 667
rect 754 666 757 670
rect 750 663 757 666
rect 760 666 763 670
rect 767 666 768 670
rect 760 663 768 666
rect 771 666 774 670
rect 771 663 778 666
rect 733 572 736 576
rect 729 569 736 572
rect 739 572 742 576
rect 746 572 747 576
rect 739 569 747 572
rect 750 572 753 576
rect 750 569 757 572
rect 894 540 897 544
rect 890 537 897 540
rect 900 540 903 544
rect 907 540 908 544
rect 900 537 908 540
rect 911 540 914 544
rect 911 537 918 540
rect 972 539 975 543
rect 968 536 975 539
rect 978 539 981 543
rect 985 539 986 543
rect 978 536 986 539
rect 989 539 992 543
rect 989 536 996 539
rect 1187 502 1191 507
rect 1194 502 1198 507
rect 1202 502 1204 507
rect 951 445 954 449
rect 947 442 954 445
rect 957 445 960 449
rect 964 445 965 449
rect 957 442 965 445
rect 968 445 971 449
rect 968 442 975 445
rect 689 391 692 395
rect 685 388 692 391
rect 695 391 698 395
rect 702 391 703 395
rect 695 388 703 391
rect 706 391 709 395
rect 706 388 713 391
rect 767 390 770 394
rect 763 387 770 390
rect 773 390 776 394
rect 780 390 781 394
rect 773 387 781 390
rect 784 390 787 394
rect 784 387 791 390
rect 746 296 749 300
rect 742 293 749 296
rect 752 296 755 300
rect 759 296 760 300
rect 752 293 760 296
rect 763 296 766 300
rect 763 293 770 296
rect -80 58 -76 63
rect -73 58 -69 63
rect -65 58 -63 63
rect 85 58 89 63
rect 92 58 96 63
rect 100 58 102 63
rect 262 59 266 64
rect 269 59 273 64
rect 277 59 279 64
rect 437 58 441 63
rect 444 58 448 63
rect 452 58 454 63
rect 835 13 839 18
rect 842 13 846 18
rect 850 13 852 18
rect 1083 12 1087 17
rect 1090 12 1094 17
rect 1098 12 1100 17
rect 913 4 918 5
rect 917 0 918 4
rect 920 4 926 5
rect 920 0 922 4
rect 932 4 937 5
rect 936 0 937 4
rect 939 4 945 5
rect 939 0 941 4
rect 957 4 962 5
rect 961 0 962 4
rect 964 4 970 5
rect 964 0 966 4
rect 976 4 981 5
rect 980 0 981 4
rect 983 4 989 5
rect 983 0 985 4
rect 1326 21 1330 26
rect 1333 21 1337 26
rect 1341 21 1343 26
rect 1161 3 1166 4
rect 1165 -1 1166 3
rect 1168 3 1174 4
rect 1168 -1 1170 3
rect 1180 3 1185 4
rect 1184 -1 1185 3
rect 1187 3 1193 4
rect 1187 -1 1189 3
rect 1205 3 1210 4
rect 1209 -1 1210 3
rect 1212 3 1218 4
rect 1212 -1 1214 3
rect 1224 3 1229 4
rect 1228 -1 1229 3
rect 1231 3 1237 4
rect 1231 -1 1233 3
rect 1595 26 1599 31
rect 1602 26 1606 31
rect 1610 26 1612 31
rect 1404 12 1409 13
rect 1408 8 1409 12
rect 1411 12 1417 13
rect 1411 8 1413 12
rect 1423 12 1428 13
rect 1427 8 1428 12
rect 1430 12 1436 13
rect 1430 8 1432 12
rect 1448 12 1453 13
rect 1452 8 1453 12
rect 1455 12 1461 13
rect 1455 8 1457 12
rect 1467 12 1472 13
rect 1471 8 1472 12
rect 1474 12 1480 13
rect 1474 8 1476 12
rect 1673 17 1678 18
rect 1677 13 1678 17
rect 1680 17 1686 18
rect 1680 13 1682 17
rect 1692 17 1697 18
rect 1696 13 1697 17
rect 1699 17 1705 18
rect 1699 13 1701 17
rect 1717 17 1722 18
rect 1721 13 1722 17
rect 1724 17 1730 18
rect 1724 13 1726 17
rect 1736 17 1741 18
rect 1740 13 1741 17
rect 1743 17 1749 18
rect 1743 13 1745 17
rect 137 -55 140 -51
rect -34 -60 -31 -56
rect -38 -63 -31 -60
rect -28 -60 -25 -56
rect -21 -60 -20 -56
rect -28 -63 -20 -60
rect -17 -60 -14 -56
rect -17 -63 -10 -60
rect 23 -61 27 -56
rect 30 -61 34 -56
rect 38 -61 40 -56
rect 133 -58 140 -55
rect 143 -55 146 -51
rect 150 -55 151 -51
rect 143 -58 151 -55
rect 154 -55 157 -51
rect 154 -58 161 -55
rect 194 -56 198 -51
rect 201 -56 205 -51
rect 209 -56 211 -51
rect 511 -55 514 -51
rect 330 -59 333 -55
rect 326 -62 333 -59
rect 336 -59 339 -55
rect 343 -59 344 -55
rect 336 -62 344 -59
rect 347 -59 350 -55
rect 347 -62 354 -59
rect 387 -60 391 -55
rect 394 -60 398 -55
rect 402 -60 404 -55
rect 507 -58 514 -55
rect 517 -55 520 -51
rect 524 -55 525 -51
rect 517 -58 525 -55
rect 528 -55 531 -51
rect 528 -58 535 -55
rect 568 -56 572 -51
rect 575 -56 579 -51
rect 583 -56 585 -51
rect 1169 -116 1172 -112
rect 1165 -119 1172 -116
rect 1175 -116 1178 -112
rect 1182 -116 1183 -112
rect 1175 -119 1183 -116
rect 1186 -116 1189 -112
rect 1186 -119 1193 -116
rect 1226 -117 1230 -112
rect 1233 -117 1237 -112
rect 1241 -117 1243 -112
rect 1545 -128 1548 -124
rect 1541 -131 1548 -128
rect 1551 -128 1554 -124
rect 1558 -128 1559 -124
rect 1551 -131 1559 -128
rect 1562 -128 1565 -124
rect 1562 -131 1569 -128
rect 1602 -129 1606 -124
rect 1609 -129 1613 -124
rect 1617 -129 1619 -124
rect 1389 -136 1392 -132
rect 1385 -139 1392 -136
rect 1395 -136 1398 -132
rect 1402 -136 1403 -132
rect 1395 -139 1403 -136
rect 1406 -136 1409 -132
rect 1406 -139 1413 -136
rect 1446 -137 1450 -132
rect 1453 -137 1457 -132
rect 1461 -137 1463 -132
rect 98 -199 101 -195
rect 94 -202 101 -199
rect 104 -199 107 -195
rect 111 -199 112 -195
rect 104 -202 112 -199
rect 115 -199 118 -195
rect 115 -202 122 -199
rect 155 -200 159 -195
rect 162 -200 166 -195
rect 170 -200 172 -195
rect 948 -231 951 -227
rect 944 -234 951 -231
rect 954 -231 957 -227
rect 961 -231 962 -227
rect 954 -234 962 -231
rect 965 -231 968 -227
rect 965 -234 972 -231
rect 1005 -232 1009 -227
rect 1012 -232 1016 -227
rect 1020 -232 1022 -227
rect 2099 -353 2102 -349
rect 2095 -356 2102 -353
rect 2105 -353 2108 -349
rect 2112 -353 2113 -349
rect 2105 -356 2113 -353
rect 2116 -353 2119 -349
rect 2116 -356 2123 -353
rect 2156 -354 2160 -349
rect 2163 -354 2167 -349
rect 2171 -354 2173 -349
rect 2316 -353 2319 -349
rect 2312 -356 2319 -353
rect 2322 -353 2325 -349
rect 2329 -353 2330 -349
rect 2322 -356 2330 -353
rect 2333 -353 2336 -349
rect 2333 -356 2340 -353
rect 2373 -354 2377 -349
rect 2380 -354 2384 -349
rect 2388 -354 2390 -349
rect 102 -397 105 -393
rect 98 -400 105 -397
rect 108 -397 111 -393
rect 115 -397 116 -393
rect 108 -400 116 -397
rect 119 -397 122 -393
rect 119 -400 126 -397
rect 159 -398 163 -393
rect 166 -398 170 -393
rect 174 -398 176 -393
rect 1289 -400 1292 -396
rect 1285 -403 1292 -400
rect 1295 -400 1298 -396
rect 1302 -400 1303 -396
rect 1295 -403 1303 -400
rect 1306 -400 1309 -396
rect 1306 -403 1313 -400
rect 1346 -401 1350 -396
rect 1353 -401 1357 -396
rect 1361 -401 1363 -396
rect 961 -417 964 -413
rect 957 -420 964 -417
rect 967 -417 970 -413
rect 974 -417 975 -413
rect 967 -420 975 -417
rect 978 -417 981 -413
rect 978 -420 985 -417
rect 1018 -418 1022 -413
rect 1025 -418 1029 -413
rect 1033 -418 1035 -413
rect -55 -573 -51 -568
rect -48 -573 -44 -568
rect -40 -573 -38 -568
rect 110 -573 114 -568
rect 117 -573 121 -568
rect 125 -573 127 -568
rect 287 -572 291 -567
rect 294 -572 298 -567
rect 302 -572 304 -567
rect 462 -573 466 -568
rect 469 -573 473 -568
rect 477 -573 479 -568
rect 162 -686 165 -682
rect -9 -691 -6 -687
rect -13 -694 -6 -691
rect -3 -691 0 -687
rect 4 -691 5 -687
rect -3 -694 5 -691
rect 8 -691 11 -687
rect 8 -694 15 -691
rect 48 -692 52 -687
rect 55 -692 59 -687
rect 63 -692 65 -687
rect 158 -689 165 -686
rect 168 -686 171 -682
rect 175 -686 176 -682
rect 168 -689 176 -686
rect 179 -686 182 -682
rect 179 -689 186 -686
rect 219 -687 223 -682
rect 226 -687 230 -682
rect 234 -687 236 -682
rect 536 -686 539 -682
rect 355 -690 358 -686
rect 351 -693 358 -690
rect 361 -690 364 -686
rect 368 -690 369 -686
rect 361 -693 369 -690
rect 372 -690 375 -686
rect 372 -693 379 -690
rect 412 -691 416 -686
rect 419 -691 423 -686
rect 427 -691 429 -686
rect 532 -689 539 -686
rect 542 -686 545 -682
rect 549 -686 550 -682
rect 542 -689 550 -686
rect 553 -686 556 -682
rect 553 -689 560 -686
rect 593 -687 597 -682
rect 600 -687 604 -682
rect 608 -687 610 -682
rect 748 -887 751 -883
rect 744 -890 751 -887
rect 754 -887 757 -883
rect 761 -887 762 -883
rect 754 -890 762 -887
rect 765 -887 768 -883
rect 765 -890 772 -887
rect 826 -888 829 -884
rect 822 -891 829 -888
rect 832 -888 835 -884
rect 839 -888 840 -884
rect 832 -891 840 -888
rect 843 -888 846 -884
rect 843 -891 850 -888
rect 805 -982 808 -978
rect 801 -985 808 -982
rect 811 -982 814 -978
rect 818 -982 819 -978
rect 811 -985 819 -982
rect 822 -982 825 -978
rect 822 -985 829 -982
rect 1649 -985 1653 -980
rect 1656 -985 1660 -980
rect 1664 -985 1666 -980
rect 1093 -997 1096 -993
rect 1089 -1000 1096 -997
rect 1099 -997 1102 -993
rect 1106 -997 1107 -993
rect 1099 -1000 1107 -997
rect 1110 -997 1113 -993
rect 1110 -1000 1117 -997
rect 1171 -998 1174 -994
rect 1167 -1001 1174 -998
rect 1177 -998 1180 -994
rect 1184 -998 1185 -994
rect 1177 -1001 1185 -998
rect 1188 -998 1191 -994
rect 1188 -1001 1195 -998
rect 1150 -1092 1153 -1088
rect 1146 -1095 1153 -1092
rect 1156 -1092 1159 -1088
rect 1163 -1092 1164 -1088
rect 1156 -1095 1164 -1092
rect 1167 -1092 1170 -1088
rect 1167 -1095 1174 -1092
rect 758 -1131 761 -1127
rect 754 -1134 761 -1131
rect 764 -1131 767 -1127
rect 771 -1131 772 -1127
rect 764 -1134 772 -1131
rect 775 -1131 778 -1127
rect 775 -1134 782 -1131
rect 836 -1132 839 -1128
rect 832 -1135 839 -1132
rect 842 -1132 845 -1128
rect 849 -1132 850 -1128
rect 842 -1135 850 -1132
rect 853 -1132 856 -1128
rect 853 -1135 860 -1132
rect 815 -1226 818 -1222
rect 811 -1229 818 -1226
rect 821 -1226 824 -1222
rect 828 -1226 829 -1222
rect 821 -1229 829 -1226
rect 832 -1226 835 -1222
rect 832 -1229 839 -1226
<< highvoltpdiffusion >>
rect 416 -79 421 -75
<< metal1 >>
rect 682 681 687 682
rect 672 680 765 681
rect 672 677 778 680
rect 672 671 676 677
rect 696 671 700 677
rect 750 676 778 677
rect 750 670 754 676
rect 774 670 778 676
rect 685 660 689 667
rect 668 656 678 660
rect 685 657 700 660
rect 763 659 767 666
rect 671 652 674 656
rect 696 654 700 657
rect 748 655 756 659
rect 763 656 778 659
rect 671 648 689 652
rect 696 651 701 654
rect 748 651 752 655
rect 774 653 778 656
rect 774 651 779 653
rect 696 647 708 651
rect 748 647 767 651
rect 774 648 786 651
rect 696 640 700 647
rect 673 627 677 636
rect 673 624 702 627
rect 682 622 689 624
rect 705 557 708 647
rect 774 639 778 648
rect 751 626 755 635
rect 751 623 780 626
rect 762 621 768 623
rect 783 597 786 648
rect 711 594 786 597
rect 711 565 715 594
rect 739 586 746 589
rect 729 582 757 586
rect 729 576 733 582
rect 753 576 757 582
rect 742 565 746 572
rect 711 561 735 565
rect 742 562 757 565
rect 753 559 757 562
rect 705 553 746 557
rect 753 555 759 559
rect 753 545 757 555
rect 900 554 905 555
rect 890 553 983 554
rect 890 550 996 553
rect 890 544 894 550
rect 914 544 918 550
rect 730 532 734 541
rect 968 549 996 550
rect 968 543 972 549
rect 992 543 996 549
rect 903 533 907 540
rect 730 529 759 532
rect 866 529 896 533
rect 903 530 918 533
rect 981 532 985 539
rect 741 527 749 529
rect 695 405 700 406
rect 685 404 778 405
rect 685 401 791 404
rect 685 395 689 401
rect 709 395 713 401
rect 763 400 791 401
rect 763 394 767 400
rect 787 394 791 400
rect 698 384 702 391
rect 681 380 691 384
rect 698 381 713 384
rect 776 383 780 390
rect 684 376 687 380
rect 709 378 713 381
rect 761 379 769 383
rect 776 380 791 383
rect 684 372 702 376
rect 709 375 714 378
rect 761 375 765 379
rect 787 377 791 380
rect 787 375 792 377
rect 709 371 721 375
rect 761 371 780 375
rect 787 372 799 375
rect 709 364 713 371
rect 686 351 690 360
rect 686 348 715 351
rect 695 346 702 348
rect 718 281 721 371
rect 787 363 791 372
rect 764 350 768 359
rect 764 347 793 350
rect 775 345 781 347
rect 796 321 799 372
rect 724 318 799 321
rect 724 289 728 318
rect 752 310 759 313
rect 742 306 770 310
rect 742 300 746 306
rect 766 300 770 306
rect 755 289 759 296
rect 724 285 748 289
rect 755 286 770 289
rect 766 283 770 286
rect 866 283 870 529
rect 889 525 892 529
rect 914 527 918 530
rect 966 528 974 532
rect 981 529 996 532
rect 889 521 907 525
rect 914 524 919 527
rect 966 524 970 528
rect 992 526 996 529
rect 992 524 997 526
rect 914 520 926 524
rect 966 520 985 524
rect 992 521 1004 524
rect 914 513 918 520
rect 891 500 895 509
rect 891 497 920 500
rect 900 495 907 497
rect 923 430 926 520
rect 992 512 996 521
rect 969 499 973 508
rect 969 496 998 499
rect 980 494 986 496
rect 1001 470 1004 521
rect 1173 513 1186 517
rect 1190 513 1214 517
rect 1183 507 1186 513
rect 1199 487 1202 502
rect 929 467 1004 470
rect 1085 483 1190 487
rect 1199 484 1988 487
rect 929 438 933 467
rect 957 459 964 462
rect 947 455 975 459
rect 947 449 951 455
rect 971 449 975 455
rect 960 438 964 445
rect 929 434 953 438
rect 960 435 975 438
rect 971 432 975 435
rect 1085 432 1089 483
rect 1199 468 1202 484
rect 1183 456 1187 463
rect 1173 450 1215 456
rect 923 426 964 430
rect 971 428 1089 432
rect 971 418 975 428
rect 948 405 952 414
rect 948 402 977 405
rect 959 400 967 402
rect 718 277 759 281
rect 766 279 870 283
rect 766 269 770 279
rect 743 256 747 265
rect 743 253 772 256
rect 754 251 762 253
rect -127 134 1813 137
rect -127 -213 -124 134
rect -94 69 -81 73
rect -77 69 -53 73
rect 71 69 84 73
rect 88 69 112 73
rect 248 70 261 74
rect 265 70 289 74
rect -84 63 -81 69
rect 81 63 84 69
rect 258 64 261 70
rect 423 69 436 73
rect 440 69 464 73
rect -68 43 -65 58
rect 97 43 100 58
rect 274 44 277 59
rect 433 63 436 69
rect -79 39 -77 43
rect -68 40 -47 43
rect -68 24 -65 40
rect -84 12 -80 19
rect -94 6 -57 12
rect -50 -67 -47 40
rect 86 39 88 43
rect 97 40 124 43
rect 263 40 265 44
rect 274 41 317 44
rect 449 43 452 58
rect 97 24 100 40
rect 81 12 85 19
rect 71 6 113 12
rect -28 -46 -23 -45
rect -38 -50 22 -46
rect 26 -50 51 -46
rect -38 -56 -34 -50
rect -14 -56 -10 -50
rect 19 -56 22 -50
rect -25 -67 -21 -60
rect -50 -71 -32 -67
rect -25 -70 -10 -67
rect -14 -73 -10 -70
rect -41 -79 -21 -75
rect -14 -76 -9 -73
rect 35 -76 38 -61
rect 121 -62 124 40
rect 274 25 277 41
rect 258 13 262 20
rect 248 7 290 13
rect 143 -41 148 -40
rect 133 -45 193 -41
rect 197 -45 222 -41
rect 133 -51 137 -45
rect 157 -51 161 -45
rect 190 -51 193 -45
rect 146 -62 150 -55
rect 121 -66 139 -62
rect 146 -65 161 -62
rect 157 -68 161 -65
rect 130 -74 150 -70
rect 157 -71 162 -68
rect 206 -70 209 -56
rect 314 -66 317 41
rect 438 39 440 43
rect 449 40 498 43
rect 1673 41 1713 45
rect 449 24 452 40
rect 433 12 437 19
rect 423 6 465 12
rect 336 -45 341 -44
rect 326 -49 386 -45
rect 390 -49 415 -45
rect 326 -55 330 -49
rect 350 -55 354 -49
rect 383 -55 386 -49
rect 339 -66 343 -59
rect 314 -70 332 -66
rect 339 -69 354 -66
rect 157 -75 197 -71
rect 206 -74 210 -70
rect 350 -72 354 -69
rect -14 -80 26 -76
rect 35 -79 54 -76
rect -14 -87 -10 -80
rect -37 -100 -33 -91
rect 35 -95 38 -79
rect -37 -103 9 -100
rect 19 -103 23 -100
rect -9 -106 23 -103
rect 51 -206 54 -79
rect 157 -82 161 -75
rect 134 -95 138 -86
rect 206 -90 209 -74
rect 323 -78 343 -74
rect 350 -75 355 -72
rect 399 -75 402 -60
rect 495 -62 498 40
rect 1404 36 1444 40
rect 1581 37 1594 41
rect 1598 37 1622 41
rect 1312 32 1325 36
rect 1329 32 1353 36
rect 913 28 953 32
rect 821 24 834 28
rect 838 24 862 28
rect 831 18 834 24
rect 847 -1 850 13
rect 913 4 917 28
rect 837 -6 838 -2
rect 847 -4 880 -1
rect 847 -21 850 -4
rect 831 -33 835 -26
rect 821 -39 863 -33
rect 517 -41 522 -40
rect 507 -45 567 -41
rect 571 -45 596 -41
rect 507 -51 511 -45
rect 531 -51 535 -45
rect 564 -51 567 -45
rect 520 -62 524 -55
rect 495 -66 513 -62
rect 520 -65 535 -62
rect 531 -68 535 -65
rect 504 -74 524 -70
rect 531 -71 536 -68
rect 580 -70 583 -56
rect 531 -75 571 -71
rect 580 -74 584 -70
rect 350 -79 390 -75
rect 399 -79 411 -75
rect 350 -86 354 -79
rect 134 -98 180 -95
rect 190 -98 194 -95
rect 162 -101 194 -98
rect 327 -99 331 -90
rect 399 -94 402 -79
rect 531 -82 535 -75
rect 508 -95 512 -86
rect 580 -90 583 -74
rect 508 -98 554 -95
rect 564 -98 568 -95
rect 327 -102 373 -99
rect 383 -102 387 -99
rect 536 -101 568 -98
rect 355 -105 387 -102
rect 877 -134 880 -4
rect 913 -27 917 0
rect 922 21 925 25
rect 929 21 945 25
rect 922 4 926 21
rect 941 4 945 21
rect 922 -27 926 0
rect 932 -27 936 0
rect 941 -27 945 0
rect 949 -12 953 28
rect 1161 27 1201 31
rect 1069 23 1082 27
rect 1086 23 1110 27
rect 957 16 980 20
rect 957 4 961 16
rect 976 4 980 16
rect 1079 17 1082 23
rect 949 -16 959 -12
rect 966 -20 970 0
rect 949 -24 970 -20
rect 932 -34 936 -31
rect 949 -34 953 -24
rect 966 -27 970 -24
rect 985 -12 989 0
rect 1095 -3 1098 12
rect 1161 3 1165 27
rect 1085 -7 1086 -3
rect 1095 -7 1097 -3
rect 985 -16 988 -12
rect 985 -27 989 -16
rect 1095 -22 1098 -7
rect 932 -38 953 -34
rect 957 -34 961 -31
rect 976 -34 980 -31
rect 1079 -34 1083 -27
rect 1161 -28 1165 -1
rect 1170 20 1173 24
rect 1177 20 1193 24
rect 1170 3 1174 20
rect 1189 3 1193 20
rect 1170 -28 1174 -1
rect 1180 -28 1184 -1
rect 1189 -28 1193 -1
rect 1197 -13 1201 27
rect 1322 26 1325 32
rect 1205 15 1228 19
rect 1205 3 1209 15
rect 1224 3 1228 15
rect 1328 2 1329 6
rect 1338 5 1341 21
rect 1404 12 1408 36
rect 1338 2 1381 5
rect 1197 -17 1207 -13
rect 1214 -21 1218 -1
rect 1197 -25 1218 -21
rect 957 -38 980 -34
rect 1069 -40 1111 -34
rect 1180 -35 1184 -32
rect 1197 -35 1201 -25
rect 1214 -28 1218 -25
rect 1233 -13 1237 -1
rect 1338 -13 1341 2
rect 1233 -17 1236 -13
rect 1233 -28 1237 -17
rect 1322 -25 1326 -18
rect 1180 -39 1201 -35
rect 1312 -31 1354 -25
rect 1205 -35 1209 -32
rect 1224 -35 1228 -32
rect 1205 -39 1228 -35
rect 1378 -93 1381 2
rect 1404 -19 1408 8
rect 1413 29 1416 33
rect 1420 29 1436 33
rect 1413 12 1417 29
rect 1432 12 1436 29
rect 1413 -19 1417 8
rect 1423 -19 1427 8
rect 1432 -19 1436 8
rect 1440 -4 1444 36
rect 1591 31 1594 37
rect 1448 24 1471 28
rect 1448 12 1452 24
rect 1467 12 1471 24
rect 1440 -8 1450 -4
rect 1457 -12 1461 8
rect 1440 -16 1461 -12
rect 1423 -26 1427 -23
rect 1440 -26 1444 -16
rect 1457 -19 1461 -16
rect 1476 -4 1480 8
rect 1597 7 1598 11
rect 1476 -8 1479 -4
rect 1607 -8 1610 26
rect 1476 -19 1480 -8
rect 1423 -30 1444 -26
rect 1673 17 1677 41
rect 1591 -20 1595 -13
rect 1673 -14 1677 13
rect 1682 34 1685 38
rect 1689 34 1705 38
rect 1682 17 1686 34
rect 1701 17 1705 34
rect 1682 -14 1686 13
rect 1692 -14 1696 13
rect 1701 -14 1705 13
rect 1709 1 1713 41
rect 1717 29 1740 33
rect 1717 17 1721 29
rect 1736 17 1740 29
rect 1709 -3 1719 1
rect 1726 -7 1730 13
rect 1709 -11 1730 -7
rect 1448 -26 1452 -23
rect 1467 -26 1471 -23
rect 1581 -26 1623 -20
rect 1692 -21 1696 -18
rect 1709 -21 1713 -11
rect 1726 -14 1730 -11
rect 1745 1 1749 13
rect 1745 -3 1748 1
rect 1745 -14 1749 -3
rect 1692 -25 1713 -21
rect 1717 -21 1721 -18
rect 1736 -21 1740 -18
rect 1717 -25 1740 -21
rect 1448 -30 1471 -26
rect 1378 -96 1524 -93
rect 1175 -102 1180 -101
rect 1165 -106 1225 -102
rect 1229 -106 1254 -102
rect 1165 -112 1169 -106
rect 1189 -112 1193 -106
rect 1222 -112 1225 -106
rect 1178 -123 1182 -116
rect 1161 -127 1171 -124
rect 1178 -126 1193 -123
rect 1189 -129 1193 -126
rect 1172 -132 1182 -131
rect 1149 -134 1182 -132
rect 877 -135 1182 -134
rect 1189 -132 1194 -129
rect 1238 -132 1241 -117
rect 1329 -114 1514 -111
rect 1329 -132 1332 -114
rect 1395 -122 1400 -121
rect 1385 -126 1445 -122
rect 1449 -126 1474 -122
rect 1385 -132 1389 -126
rect 1409 -132 1413 -126
rect 877 -137 1155 -135
rect 1189 -136 1229 -132
rect 1238 -135 1338 -132
rect 104 -185 109 -184
rect 94 -189 154 -185
rect 158 -189 183 -185
rect 94 -195 98 -189
rect 118 -195 122 -189
rect 151 -195 154 -189
rect 107 -206 111 -199
rect 51 -210 100 -206
rect 107 -209 122 -206
rect 118 -212 122 -209
rect -127 -214 102 -213
rect -127 -218 111 -214
rect 118 -215 123 -212
rect 167 -214 170 -200
rect 64 -405 69 -218
rect 118 -219 158 -215
rect 167 -218 172 -214
rect 118 -226 122 -219
rect 95 -239 99 -230
rect 167 -234 170 -218
rect 95 -242 141 -239
rect 151 -242 155 -239
rect 123 -245 155 -242
rect 877 -247 880 -137
rect 1189 -143 1193 -136
rect 1166 -156 1170 -147
rect 1238 -151 1241 -135
rect 1166 -159 1212 -156
rect 1222 -159 1226 -156
rect 1194 -162 1226 -159
rect 954 -217 959 -216
rect 944 -221 1004 -217
rect 1008 -221 1033 -217
rect 944 -227 948 -221
rect 968 -227 972 -221
rect 1001 -227 1004 -221
rect 957 -238 961 -231
rect 940 -242 950 -239
rect 957 -241 972 -238
rect 968 -244 972 -241
rect 951 -247 961 -246
rect 877 -250 961 -247
rect 968 -247 973 -244
rect 1017 -246 1020 -232
rect 108 -383 113 -382
rect 98 -387 158 -383
rect 162 -387 187 -383
rect 98 -393 102 -387
rect 122 -393 126 -387
rect 155 -393 158 -387
rect 111 -404 115 -397
rect 64 -408 104 -405
rect 111 -407 126 -404
rect 122 -410 126 -407
rect 105 -413 115 -412
rect 82 -416 115 -413
rect 122 -413 127 -410
rect 171 -412 174 -398
rect -69 -562 -56 -558
rect -52 -562 -28 -558
rect -59 -568 -56 -562
rect -43 -588 -40 -573
rect -54 -592 -52 -588
rect -43 -591 -22 -588
rect -43 -607 -40 -591
rect -59 -619 -55 -612
rect -69 -625 -32 -619
rect -25 -698 -22 -591
rect -3 -677 2 -676
rect -13 -681 47 -677
rect 51 -681 76 -677
rect -13 -687 -9 -681
rect 11 -687 15 -681
rect 44 -687 47 -681
rect 0 -698 4 -691
rect -25 -702 -7 -698
rect 0 -701 15 -698
rect 11 -704 15 -701
rect -16 -710 4 -706
rect 11 -707 16 -704
rect 60 -707 63 -692
rect 82 -707 85 -416
rect 122 -417 162 -413
rect 171 -416 176 -412
rect 122 -424 126 -417
rect 99 -437 103 -428
rect 171 -432 174 -416
rect 877 -425 880 -250
rect 968 -251 1008 -247
rect 1017 -250 1021 -246
rect 968 -258 972 -251
rect 945 -271 949 -262
rect 1017 -266 1020 -250
rect 945 -274 991 -271
rect 1001 -274 1005 -271
rect 973 -277 1005 -274
rect 967 -403 972 -402
rect 957 -407 1017 -403
rect 1021 -407 1046 -403
rect 957 -413 961 -407
rect 981 -413 985 -407
rect 1014 -413 1017 -407
rect 1257 -408 1260 -135
rect 1335 -152 1338 -135
rect 1442 -132 1445 -126
rect 1398 -143 1402 -136
rect 1381 -147 1391 -144
rect 1398 -146 1413 -143
rect 1409 -149 1413 -146
rect 1392 -152 1402 -151
rect 1335 -155 1402 -152
rect 1409 -152 1414 -149
rect 1458 -151 1461 -137
rect 1511 -144 1514 -114
rect 1521 -136 1524 -96
rect 1551 -114 1556 -113
rect 1541 -118 1601 -114
rect 1605 -118 1630 -114
rect 1541 -124 1545 -118
rect 1565 -124 1569 -118
rect 1598 -124 1601 -118
rect 1554 -135 1558 -128
rect 1521 -139 1547 -136
rect 1554 -138 1569 -135
rect 1565 -141 1569 -138
rect 1548 -144 1558 -143
rect 1511 -147 1558 -144
rect 1565 -144 1570 -141
rect 1614 -144 1617 -129
rect 1810 -144 1813 134
rect 1565 -148 1605 -144
rect 1614 -147 1813 -144
rect 1409 -156 1449 -152
rect 1458 -155 1463 -151
rect 1565 -155 1569 -148
rect 1409 -163 1413 -156
rect 1386 -176 1390 -167
rect 1458 -171 1461 -155
rect 1542 -168 1546 -159
rect 1614 -163 1617 -147
rect 1542 -171 1588 -168
rect 1598 -171 1602 -168
rect 1570 -174 1602 -171
rect 1386 -179 1432 -176
rect 1442 -179 1446 -176
rect 1414 -182 1446 -179
rect 1985 -361 1988 484
rect 2105 -339 2110 -338
rect 2322 -339 2327 -338
rect 2095 -343 2155 -339
rect 2159 -343 2184 -339
rect 2312 -343 2372 -339
rect 2376 -343 2401 -339
rect 2095 -349 2099 -343
rect 2119 -349 2123 -343
rect 2152 -349 2155 -343
rect 2312 -349 2316 -343
rect 2336 -349 2340 -343
rect 2108 -360 2112 -353
rect 2369 -349 2372 -343
rect 1985 -364 2101 -361
rect 2108 -363 2123 -360
rect 2119 -366 2123 -363
rect 2102 -369 2112 -368
rect 1984 -372 2112 -369
rect 2119 -369 2124 -366
rect 2168 -369 2171 -354
rect 2325 -360 2329 -353
rect 2308 -364 2318 -361
rect 2325 -363 2340 -360
rect 2336 -366 2340 -363
rect 2319 -369 2329 -368
rect 1295 -386 1300 -385
rect 1285 -390 1345 -386
rect 1349 -390 1374 -386
rect 1285 -396 1289 -390
rect 1309 -396 1313 -390
rect 1342 -396 1345 -390
rect 1298 -407 1302 -400
rect 1257 -411 1291 -408
rect 1298 -410 1313 -407
rect 1309 -413 1313 -410
rect 970 -424 974 -417
rect 1292 -416 1302 -415
rect 877 -428 963 -425
rect 970 -427 985 -424
rect 981 -430 985 -427
rect 964 -433 974 -432
rect 909 -436 974 -433
rect 981 -433 986 -430
rect 1030 -432 1033 -418
rect 1259 -419 1302 -416
rect 1309 -416 1314 -413
rect 1358 -414 1361 -401
rect 99 -440 145 -437
rect 155 -440 159 -437
rect 127 -443 159 -440
rect 96 -562 109 -558
rect 113 -562 137 -558
rect 273 -561 286 -557
rect 290 -561 314 -557
rect 106 -568 109 -562
rect 283 -567 286 -561
rect 448 -562 461 -558
rect 465 -562 489 -558
rect 122 -588 125 -573
rect 299 -587 302 -572
rect 458 -568 461 -562
rect 111 -592 113 -588
rect 122 -591 149 -588
rect 288 -591 290 -587
rect 299 -590 342 -587
rect 474 -588 477 -573
rect 122 -607 125 -591
rect 106 -619 110 -612
rect 96 -625 138 -619
rect 146 -693 149 -591
rect 299 -606 302 -590
rect 283 -618 287 -611
rect 273 -624 315 -618
rect 168 -672 173 -671
rect 158 -676 218 -672
rect 222 -676 247 -672
rect 158 -682 162 -676
rect 182 -682 186 -676
rect 215 -682 218 -676
rect 171 -693 175 -686
rect 146 -697 164 -693
rect 171 -696 186 -693
rect 182 -699 186 -696
rect 155 -705 175 -701
rect 182 -702 187 -699
rect 231 -702 234 -687
rect 339 -697 342 -590
rect 463 -592 465 -588
rect 474 -591 523 -588
rect 474 -607 477 -591
rect 458 -619 462 -612
rect 448 -625 490 -619
rect 361 -676 366 -675
rect 351 -680 411 -676
rect 415 -680 440 -676
rect 351 -686 355 -680
rect 375 -686 379 -680
rect 408 -686 411 -680
rect 364 -697 368 -690
rect 339 -701 357 -697
rect 364 -700 379 -697
rect 11 -711 51 -707
rect 60 -710 85 -707
rect 182 -706 222 -702
rect 231 -705 266 -702
rect 375 -703 379 -700
rect 11 -718 15 -711
rect -12 -731 -8 -722
rect 60 -726 63 -710
rect 182 -713 186 -706
rect 159 -726 163 -717
rect 231 -721 234 -705
rect 159 -729 205 -726
rect 215 -729 219 -726
rect -12 -734 34 -731
rect 44 -734 48 -731
rect 187 -732 219 -729
rect 16 -737 48 -734
rect 263 -795 266 -705
rect 348 -709 368 -705
rect 375 -706 380 -703
rect 424 -705 427 -691
rect 520 -693 523 -591
rect 542 -672 547 -671
rect 532 -676 592 -672
rect 596 -676 621 -672
rect 532 -682 536 -676
rect 556 -682 560 -676
rect 589 -682 592 -676
rect 545 -693 549 -686
rect 520 -697 538 -693
rect 545 -696 560 -693
rect 556 -699 560 -696
rect 529 -705 549 -701
rect 556 -702 561 -699
rect 605 -701 608 -687
rect 375 -710 415 -706
rect 424 -708 452 -705
rect 375 -717 379 -710
rect 352 -730 356 -721
rect 424 -725 427 -708
rect 352 -733 398 -730
rect 408 -733 412 -730
rect 380 -736 412 -733
rect 449 -750 452 -708
rect 556 -706 596 -702
rect 605 -705 610 -701
rect 556 -713 560 -706
rect 533 -726 537 -717
rect 605 -721 608 -705
rect 533 -729 579 -726
rect 589 -729 593 -726
rect 561 -732 593 -729
rect 909 -750 912 -436
rect 981 -437 1021 -433
rect 1030 -436 1035 -432
rect 981 -444 985 -437
rect 958 -457 962 -448
rect 1030 -452 1033 -436
rect 958 -460 1004 -457
rect 1014 -460 1018 -457
rect 986 -463 1018 -460
rect 449 -753 912 -750
rect 1259 -795 1262 -419
rect 1309 -420 1349 -416
rect 1358 -420 1364 -414
rect 1309 -427 1313 -420
rect 1286 -440 1290 -431
rect 1358 -435 1361 -420
rect 1286 -443 1332 -440
rect 1342 -443 1346 -440
rect 1314 -446 1346 -443
rect 263 -798 1262 -795
rect 754 -873 759 -872
rect 744 -874 837 -873
rect 744 -877 850 -874
rect 744 -883 748 -877
rect 768 -883 772 -877
rect 822 -878 850 -877
rect 822 -884 826 -878
rect 846 -884 850 -878
rect 757 -894 761 -887
rect 740 -898 750 -894
rect 757 -897 772 -894
rect 835 -895 839 -888
rect 743 -902 746 -898
rect 768 -900 772 -897
rect 820 -899 828 -895
rect 835 -898 850 -895
rect 743 -906 761 -902
rect 768 -903 773 -900
rect 820 -903 824 -899
rect 846 -901 850 -898
rect 846 -903 851 -901
rect 768 -907 780 -903
rect 820 -907 839 -903
rect 846 -906 858 -903
rect 768 -914 772 -907
rect 745 -927 749 -918
rect 745 -930 774 -927
rect 754 -932 761 -930
rect 777 -997 780 -907
rect 846 -915 850 -906
rect 823 -928 827 -919
rect 823 -931 852 -928
rect 834 -933 840 -931
rect 855 -957 858 -906
rect 783 -960 858 -957
rect 783 -989 787 -960
rect 811 -968 818 -965
rect 801 -972 829 -968
rect 801 -978 805 -972
rect 825 -978 829 -972
rect 1635 -974 1648 -970
rect 1652 -974 1676 -970
rect 1645 -980 1648 -974
rect 814 -989 818 -982
rect 1099 -983 1104 -982
rect 1089 -984 1182 -983
rect 1089 -987 1195 -984
rect 783 -993 807 -989
rect 814 -992 829 -989
rect 825 -995 829 -992
rect 1089 -993 1093 -987
rect 1113 -993 1117 -987
rect 777 -1001 818 -997
rect 825 -999 831 -995
rect 1167 -988 1195 -987
rect 1167 -994 1171 -988
rect 1191 -994 1195 -988
rect 825 -1009 829 -999
rect 1102 -1004 1106 -997
rect 1069 -1008 1095 -1004
rect 1102 -1007 1117 -1004
rect 1180 -1005 1184 -998
rect 1661 -1000 1664 -985
rect 1984 -1000 1988 -372
rect 2119 -373 2159 -369
rect 2168 -372 2329 -369
rect 2336 -369 2341 -366
rect 2385 -369 2388 -354
rect 2119 -380 2123 -373
rect 2096 -393 2100 -384
rect 2168 -388 2171 -372
rect 2336 -373 2376 -369
rect 2385 -372 2416 -369
rect 2336 -380 2340 -373
rect 2313 -393 2317 -384
rect 2385 -388 2388 -372
rect 2096 -396 2142 -393
rect 2152 -396 2156 -393
rect 2313 -396 2359 -393
rect 2369 -396 2373 -393
rect 2124 -399 2156 -396
rect 2341 -399 2373 -396
rect 1577 -1004 1652 -1000
rect 1661 -1004 1988 -1000
rect 802 -1022 806 -1013
rect 802 -1025 831 -1022
rect 813 -1027 821 -1025
rect 764 -1117 769 -1116
rect 754 -1118 847 -1117
rect 754 -1121 860 -1118
rect 754 -1127 758 -1121
rect 778 -1127 782 -1121
rect 832 -1122 860 -1121
rect 832 -1128 836 -1122
rect 856 -1128 860 -1122
rect 767 -1138 771 -1131
rect 750 -1142 760 -1138
rect 767 -1141 782 -1138
rect 845 -1139 849 -1132
rect 753 -1146 756 -1142
rect 778 -1144 782 -1141
rect 830 -1143 838 -1139
rect 845 -1142 860 -1139
rect 753 -1150 771 -1146
rect 778 -1147 783 -1144
rect 830 -1147 834 -1143
rect 856 -1145 860 -1142
rect 856 -1147 861 -1145
rect 778 -1151 790 -1147
rect 830 -1151 849 -1147
rect 856 -1150 868 -1147
rect 778 -1158 782 -1151
rect 755 -1171 759 -1162
rect 755 -1174 784 -1171
rect 764 -1176 771 -1174
rect 787 -1241 790 -1151
rect 856 -1159 860 -1150
rect 833 -1172 837 -1163
rect 833 -1175 862 -1172
rect 844 -1177 850 -1175
rect 865 -1201 868 -1150
rect 793 -1204 868 -1201
rect 793 -1233 797 -1204
rect 821 -1212 828 -1209
rect 811 -1216 839 -1212
rect 811 -1222 815 -1216
rect 835 -1222 839 -1216
rect 824 -1233 828 -1226
rect 793 -1237 817 -1233
rect 824 -1236 839 -1233
rect 835 -1239 839 -1236
rect 1069 -1239 1073 -1008
rect 1088 -1012 1091 -1008
rect 1113 -1010 1117 -1007
rect 1165 -1009 1173 -1005
rect 1180 -1008 1195 -1005
rect 1088 -1016 1106 -1012
rect 1113 -1013 1118 -1010
rect 1165 -1013 1169 -1009
rect 1191 -1011 1195 -1008
rect 1191 -1013 1196 -1011
rect 1113 -1017 1125 -1013
rect 1165 -1017 1184 -1013
rect 1191 -1016 1203 -1013
rect 1113 -1024 1117 -1017
rect 1090 -1037 1094 -1028
rect 1090 -1040 1119 -1037
rect 1099 -1042 1106 -1040
rect 1122 -1107 1125 -1017
rect 1191 -1025 1195 -1016
rect 1168 -1038 1172 -1029
rect 1168 -1041 1197 -1038
rect 1179 -1043 1185 -1041
rect 1200 -1067 1203 -1016
rect 1128 -1070 1203 -1067
rect 1128 -1099 1132 -1070
rect 1156 -1078 1163 -1075
rect 1146 -1082 1174 -1078
rect 1146 -1088 1150 -1082
rect 1170 -1088 1174 -1082
rect 1159 -1099 1163 -1092
rect 1128 -1103 1152 -1099
rect 1159 -1102 1174 -1099
rect 1170 -1105 1174 -1102
rect 1577 -1105 1581 -1004
rect 1661 -1019 1664 -1004
rect 1645 -1031 1649 -1024
rect 1635 -1037 1677 -1031
rect 1122 -1111 1163 -1107
rect 1170 -1109 1581 -1105
rect 1170 -1119 1174 -1109
rect 1147 -1132 1151 -1123
rect 1147 -1135 1176 -1132
rect 1158 -1137 1166 -1135
rect 787 -1245 828 -1241
rect 835 -1243 1073 -1239
rect 835 -1253 839 -1243
rect 812 -1266 816 -1257
rect 812 -1269 841 -1266
rect 823 -1271 831 -1269
<< metal2 >>
rect -170 656 662 660
rect -170 -278 -166 656
rect 733 654 741 659
rect 733 606 737 654
rect 733 602 1509 606
rect 837 564 945 569
rect 837 559 842 564
rect 763 555 842 559
rect 762 554 842 555
rect 940 532 945 564
rect 940 527 959 532
rect 620 380 675 384
rect 620 -70 624 380
rect 746 378 754 383
rect 746 330 750 378
rect 746 326 1042 330
rect 810 40 929 43
rect 810 -2 814 40
rect 925 25 929 40
rect 810 -6 833 -2
rect 214 -74 233 -70
rect 588 -74 624 -70
rect 176 -218 190 -214
rect 186 -278 190 -218
rect -170 -282 190 -278
rect 229 -306 233 -74
rect 416 -79 433 -75
rect 429 -239 433 -79
rect 429 -243 936 -239
rect 1038 -246 1042 326
rect 1301 48 1420 51
rect 1058 39 1177 42
rect 1058 -3 1062 39
rect 1173 24 1177 39
rect 1301 6 1305 48
rect 1416 33 1420 48
rect 1301 2 1324 6
rect 1058 -7 1081 -3
rect 1102 -7 1143 -3
rect 1140 -124 1143 -7
rect 1140 -128 1157 -124
rect 1025 -250 1042 -246
rect 1311 -148 1377 -144
rect 1311 -306 1315 -148
rect 1505 -151 1509 602
rect 1570 53 1689 56
rect 1570 11 1574 53
rect 1685 38 1689 53
rect 1570 7 1593 11
rect 1467 -155 1509 -151
rect 229 -310 1315 -306
rect 180 -416 215 -412
rect 211 -498 215 -416
rect 1372 -420 1396 -414
rect 1039 -436 1060 -432
rect -140 -502 215 -498
rect -140 -1035 -136 -502
rect 614 -705 710 -701
rect 706 -894 710 -705
rect 706 -898 734 -894
rect 805 -900 813 -895
rect 805 -947 809 -900
rect 1056 -947 1060 -436
rect 805 -951 1060 -947
rect 855 -952 858 -951
rect 1064 -975 1156 -970
rect 1064 -995 1069 -975
rect 835 -999 1069 -995
rect 834 -1000 1069 -999
rect 1151 -1005 1156 -975
rect 1151 -1010 1158 -1005
rect -140 -1039 720 -1035
rect 716 -1138 720 -1039
rect 716 -1142 744 -1138
rect 815 -1144 823 -1139
rect 815 -1191 819 -1144
rect 1390 -1191 1396 -420
rect 815 -1195 1396 -1191
rect 865 -1196 868 -1195
<< ntransistor >>
rect 679 631 682 640
rect 690 631 693 640
rect 757 630 760 639
rect 768 630 771 639
rect 736 536 739 545
rect 747 536 750 545
rect 897 504 900 513
rect 908 504 911 513
rect 975 503 978 512
rect 986 503 989 512
rect 1191 463 1194 468
rect 954 409 957 418
rect 965 409 968 418
rect 692 355 695 364
rect 703 355 706 364
rect 770 354 773 363
rect 781 354 784 363
rect 749 260 752 269
rect 760 260 763 269
rect -76 19 -73 24
rect 89 19 92 24
rect 266 20 269 25
rect 441 19 444 24
rect 839 -26 842 -21
rect 918 -31 920 -26
rect 937 -31 939 -26
rect 962 -31 964 -26
rect 981 -31 983 -26
rect 1087 -27 1090 -22
rect 1166 -32 1168 -27
rect 1185 -32 1187 -27
rect 1210 -32 1212 -27
rect 1229 -32 1231 -27
rect 1330 -18 1333 -13
rect 1409 -23 1411 -18
rect 1428 -23 1430 -18
rect 1453 -23 1455 -18
rect 1472 -23 1474 -18
rect 1599 -13 1602 -8
rect 1678 -18 1680 -13
rect 1697 -18 1699 -13
rect 1722 -18 1724 -13
rect 1741 -18 1743 -13
rect -31 -96 -28 -87
rect -20 -96 -17 -87
rect 140 -91 143 -82
rect 151 -91 154 -82
rect 198 -95 201 -90
rect 333 -95 336 -86
rect 344 -95 347 -86
rect 514 -91 517 -82
rect 525 -91 528 -82
rect 27 -100 30 -95
rect 391 -99 394 -94
rect 572 -95 575 -90
rect 1172 -152 1175 -143
rect 1183 -152 1186 -143
rect 1230 -156 1233 -151
rect 1392 -172 1395 -163
rect 1403 -172 1406 -163
rect 1548 -164 1551 -155
rect 1559 -164 1562 -155
rect 1606 -168 1609 -163
rect 1450 -176 1453 -171
rect 101 -235 104 -226
rect 112 -235 115 -226
rect 159 -239 162 -234
rect 951 -267 954 -258
rect 962 -267 965 -258
rect 1009 -271 1012 -266
rect 2102 -389 2105 -380
rect 2113 -389 2116 -380
rect 2160 -393 2163 -388
rect 2319 -389 2322 -380
rect 2330 -389 2333 -380
rect 2377 -393 2380 -388
rect 105 -433 108 -424
rect 116 -433 119 -424
rect 163 -437 166 -432
rect 1292 -436 1295 -427
rect 1303 -436 1306 -427
rect 964 -453 967 -444
rect 975 -453 978 -444
rect 1350 -440 1353 -435
rect 1022 -457 1025 -452
rect -51 -612 -48 -607
rect 114 -612 117 -607
rect 291 -611 294 -606
rect 466 -612 469 -607
rect -6 -727 -3 -718
rect 5 -727 8 -718
rect 165 -722 168 -713
rect 176 -722 179 -713
rect 223 -726 226 -721
rect 358 -726 361 -717
rect 369 -726 372 -717
rect 539 -722 542 -713
rect 550 -722 553 -713
rect 52 -731 55 -726
rect 416 -730 419 -725
rect 597 -726 600 -721
rect 751 -923 754 -914
rect 762 -923 765 -914
rect 829 -924 832 -915
rect 840 -924 843 -915
rect 808 -1018 811 -1009
rect 819 -1018 822 -1009
rect 1096 -1033 1099 -1024
rect 1107 -1033 1110 -1024
rect 1653 -1024 1656 -1019
rect 1174 -1034 1177 -1025
rect 1185 -1034 1188 -1025
rect 1153 -1128 1156 -1119
rect 1164 -1128 1167 -1119
rect 761 -1167 764 -1158
rect 772 -1167 775 -1158
rect 839 -1168 842 -1159
rect 850 -1168 853 -1159
rect 818 -1262 821 -1253
rect 829 -1262 832 -1253
<< ptransistor >>
rect 679 664 682 671
rect 690 664 693 671
rect 757 663 760 670
rect 768 663 771 670
rect 736 569 739 576
rect 747 569 750 576
rect 897 537 900 544
rect 908 537 911 544
rect 975 536 978 543
rect 986 536 989 543
rect 1191 502 1194 507
rect 954 442 957 449
rect 965 442 968 449
rect 692 388 695 395
rect 703 388 706 395
rect 770 387 773 394
rect 781 387 784 394
rect 749 293 752 300
rect 760 293 763 300
rect -76 58 -73 63
rect 89 58 92 63
rect 266 59 269 64
rect 441 58 444 63
rect 839 13 842 18
rect 1087 12 1090 17
rect 918 0 920 5
rect 937 0 939 5
rect 962 0 964 5
rect 981 0 983 5
rect 1330 21 1333 26
rect 1166 -1 1168 4
rect 1185 -1 1187 4
rect 1210 -1 1212 4
rect 1229 -1 1231 4
rect 1599 26 1602 31
rect 1409 8 1411 13
rect 1428 8 1430 13
rect 1453 8 1455 13
rect 1472 8 1474 13
rect 1678 13 1680 18
rect 1697 13 1699 18
rect 1722 13 1724 18
rect 1741 13 1743 18
rect -31 -63 -28 -56
rect -20 -63 -17 -56
rect 27 -61 30 -56
rect 140 -58 143 -51
rect 151 -58 154 -51
rect 198 -56 201 -51
rect 333 -62 336 -55
rect 344 -62 347 -55
rect 391 -60 394 -55
rect 514 -58 517 -51
rect 525 -58 528 -51
rect 572 -56 575 -51
rect 1172 -119 1175 -112
rect 1183 -119 1186 -112
rect 1230 -117 1233 -112
rect 1548 -131 1551 -124
rect 1559 -131 1562 -124
rect 1606 -129 1609 -124
rect 1392 -139 1395 -132
rect 1403 -139 1406 -132
rect 1450 -137 1453 -132
rect 101 -202 104 -195
rect 112 -202 115 -195
rect 159 -200 162 -195
rect 951 -234 954 -227
rect 962 -234 965 -227
rect 1009 -232 1012 -227
rect 2102 -356 2105 -349
rect 2113 -356 2116 -349
rect 2160 -354 2163 -349
rect 2319 -356 2322 -349
rect 2330 -356 2333 -349
rect 2377 -354 2380 -349
rect 105 -400 108 -393
rect 116 -400 119 -393
rect 163 -398 166 -393
rect 1292 -403 1295 -396
rect 1303 -403 1306 -396
rect 1350 -401 1353 -396
rect 964 -420 967 -413
rect 975 -420 978 -413
rect 1022 -418 1025 -413
rect -51 -573 -48 -568
rect 114 -573 117 -568
rect 291 -572 294 -567
rect 466 -573 469 -568
rect -6 -694 -3 -687
rect 5 -694 8 -687
rect 52 -692 55 -687
rect 165 -689 168 -682
rect 176 -689 179 -682
rect 223 -687 226 -682
rect 358 -693 361 -686
rect 369 -693 372 -686
rect 416 -691 419 -686
rect 539 -689 542 -682
rect 550 -689 553 -682
rect 597 -687 600 -682
rect 751 -890 754 -883
rect 762 -890 765 -883
rect 829 -891 832 -884
rect 840 -891 843 -884
rect 808 -985 811 -978
rect 819 -985 822 -978
rect 1653 -985 1656 -980
rect 1096 -1000 1099 -993
rect 1107 -1000 1110 -993
rect 1174 -1001 1177 -994
rect 1185 -1001 1188 -994
rect 1153 -1095 1156 -1088
rect 1164 -1095 1167 -1088
rect 761 -1134 764 -1127
rect 772 -1134 775 -1127
rect 839 -1135 842 -1128
rect 850 -1135 853 -1128
rect 818 -1229 821 -1222
rect 829 -1229 832 -1222
<< polycontact >>
rect 678 656 682 660
rect 756 655 760 659
rect 689 648 693 652
rect 767 647 771 651
rect 735 561 739 565
rect 746 553 750 557
rect 896 529 900 533
rect 974 528 978 532
rect 907 521 911 525
rect 985 520 989 524
rect 1190 483 1194 487
rect 953 434 957 438
rect 964 426 968 430
rect 691 380 695 384
rect 769 379 773 383
rect 702 372 706 376
rect 780 371 784 375
rect 748 285 752 289
rect 759 277 763 281
rect -77 39 -73 43
rect 88 39 92 43
rect 265 40 269 44
rect 440 39 444 43
rect 838 -6 842 -2
rect 959 -16 963 -12
rect 1086 -7 1090 -3
rect 988 -16 992 -12
rect 1329 2 1333 6
rect 1207 -17 1211 -13
rect 1236 -17 1240 -13
rect 1450 -8 1454 -4
rect 1598 7 1602 11
rect 1479 -8 1483 -4
rect 1719 -3 1723 1
rect 1748 -3 1752 1
rect -32 -71 -28 -67
rect -21 -79 -17 -75
rect 139 -66 143 -62
rect 26 -80 30 -76
rect 150 -74 154 -70
rect 332 -70 336 -66
rect 197 -75 201 -71
rect 343 -78 347 -74
rect 513 -66 517 -62
rect 390 -79 394 -75
rect 524 -74 528 -70
rect 571 -75 575 -71
rect 1171 -127 1175 -123
rect 1182 -135 1186 -131
rect 1229 -136 1233 -132
rect 1391 -147 1395 -143
rect 1402 -155 1406 -151
rect 1547 -139 1551 -135
rect 1449 -156 1453 -152
rect 1558 -147 1562 -143
rect 1605 -148 1609 -144
rect 100 -210 104 -206
rect 111 -218 115 -214
rect 158 -219 162 -215
rect 950 -242 954 -238
rect 961 -250 965 -246
rect 1008 -251 1012 -247
rect 2101 -364 2105 -360
rect 2112 -372 2116 -368
rect 2318 -364 2322 -360
rect 2159 -373 2163 -369
rect 2329 -372 2333 -368
rect 2376 -373 2380 -369
rect 104 -408 108 -404
rect 115 -416 119 -412
rect 1291 -411 1295 -407
rect 162 -417 166 -413
rect 963 -428 967 -424
rect 974 -436 978 -432
rect 1302 -419 1306 -415
rect 1349 -420 1353 -416
rect 1021 -437 1025 -433
rect -52 -592 -48 -588
rect 113 -592 117 -588
rect 290 -591 294 -587
rect 465 -592 469 -588
rect -7 -702 -3 -698
rect 4 -710 8 -706
rect 164 -697 168 -693
rect 51 -711 55 -707
rect 175 -705 179 -701
rect 357 -701 361 -697
rect 222 -706 226 -702
rect 368 -709 372 -705
rect 538 -697 542 -693
rect 415 -710 419 -706
rect 549 -705 553 -701
rect 596 -706 600 -702
rect 750 -898 754 -894
rect 828 -899 832 -895
rect 761 -906 765 -902
rect 839 -907 843 -903
rect 807 -993 811 -989
rect 818 -1001 822 -997
rect 1095 -1008 1099 -1004
rect 1173 -1009 1177 -1005
rect 1106 -1016 1110 -1012
rect 1652 -1004 1656 -1000
rect 1184 -1017 1188 -1013
rect 1152 -1103 1156 -1099
rect 1163 -1111 1167 -1107
rect 760 -1142 764 -1138
rect 838 -1143 842 -1139
rect 771 -1150 775 -1146
rect 849 -1151 853 -1147
rect 817 -1237 821 -1233
rect 828 -1245 832 -1241
<< ndcontact >>
rect 673 636 677 640
rect 696 636 700 640
rect 751 635 755 639
rect 774 635 778 639
rect 730 541 734 545
rect 753 541 757 545
rect 891 509 895 513
rect 914 509 918 513
rect 969 508 973 512
rect 992 508 996 512
rect 1183 463 1188 468
rect 1198 463 1202 468
rect 948 414 952 418
rect 971 414 975 418
rect 686 360 690 364
rect 709 360 713 364
rect 764 359 768 363
rect 787 359 791 363
rect 743 265 747 269
rect 766 265 770 269
rect -84 19 -79 24
rect -69 19 -65 24
rect 81 19 86 24
rect 96 19 100 24
rect 258 20 263 25
rect 273 20 277 25
rect 433 19 438 24
rect 448 19 452 24
rect 831 -26 836 -21
rect 846 -26 850 -21
rect 913 -31 917 -27
rect 922 -31 926 -27
rect 932 -31 936 -27
rect 941 -31 945 -27
rect 957 -31 961 -27
rect 966 -31 970 -27
rect 976 -31 980 -27
rect 985 -31 989 -27
rect 1079 -27 1084 -22
rect 1094 -27 1098 -22
rect 1161 -32 1165 -28
rect 1170 -32 1174 -28
rect 1180 -32 1184 -28
rect 1189 -32 1193 -28
rect 1205 -32 1209 -28
rect 1214 -32 1218 -28
rect 1224 -32 1228 -28
rect 1233 -32 1237 -28
rect 1322 -18 1327 -13
rect 1337 -18 1341 -13
rect 1404 -23 1408 -19
rect 1413 -23 1417 -19
rect 1423 -23 1427 -19
rect 1432 -23 1436 -19
rect 1448 -23 1452 -19
rect 1457 -23 1461 -19
rect 1467 -23 1471 -19
rect 1476 -23 1480 -19
rect 1591 -13 1596 -8
rect 1606 -13 1610 -8
rect 1673 -18 1677 -14
rect 1682 -18 1686 -14
rect 1692 -18 1696 -14
rect 1701 -18 1705 -14
rect 1717 -18 1721 -14
rect 1726 -18 1730 -14
rect 1736 -18 1740 -14
rect 1745 -18 1749 -14
rect -37 -91 -33 -87
rect -14 -91 -10 -87
rect 134 -86 138 -82
rect 157 -86 161 -82
rect 327 -90 331 -86
rect 190 -95 195 -90
rect 205 -95 209 -90
rect 350 -90 354 -86
rect 508 -86 512 -82
rect 531 -86 535 -82
rect 19 -100 24 -95
rect 34 -100 38 -95
rect 383 -99 388 -94
rect 398 -99 402 -94
rect 564 -95 569 -90
rect 579 -95 583 -90
rect 1166 -147 1170 -143
rect 1189 -147 1193 -143
rect 1222 -156 1227 -151
rect 1237 -156 1241 -151
rect 1386 -167 1390 -163
rect 1409 -167 1413 -163
rect 1542 -159 1546 -155
rect 1565 -159 1569 -155
rect 1598 -168 1603 -163
rect 1613 -168 1617 -163
rect 1442 -176 1447 -171
rect 1457 -176 1461 -171
rect 95 -230 99 -226
rect 118 -230 122 -226
rect 151 -239 156 -234
rect 166 -239 170 -234
rect 945 -262 949 -258
rect 968 -262 972 -258
rect 1001 -271 1006 -266
rect 1016 -271 1020 -266
rect 2096 -384 2100 -380
rect 2119 -384 2123 -380
rect 2313 -384 2317 -380
rect 2152 -393 2157 -388
rect 2167 -393 2171 -388
rect 2336 -384 2340 -380
rect 2369 -393 2374 -388
rect 2384 -393 2388 -388
rect 99 -428 103 -424
rect 122 -428 126 -424
rect 155 -437 160 -432
rect 170 -437 174 -432
rect 1286 -431 1290 -427
rect 1309 -431 1313 -427
rect 958 -448 962 -444
rect 981 -448 985 -444
rect 1342 -440 1347 -435
rect 1357 -440 1361 -435
rect 1014 -457 1019 -452
rect 1029 -457 1033 -452
rect -59 -612 -54 -607
rect -44 -612 -40 -607
rect 106 -612 111 -607
rect 121 -612 125 -607
rect 283 -611 288 -606
rect 298 -611 302 -606
rect 458 -612 463 -607
rect 473 -612 477 -607
rect -12 -722 -8 -718
rect 11 -722 15 -718
rect 159 -717 163 -713
rect 182 -717 186 -713
rect 352 -721 356 -717
rect 215 -726 220 -721
rect 230 -726 234 -721
rect 375 -721 379 -717
rect 533 -717 537 -713
rect 556 -717 560 -713
rect 44 -731 49 -726
rect 59 -731 63 -726
rect 408 -730 413 -725
rect 423 -730 427 -725
rect 589 -726 594 -721
rect 604 -726 608 -721
rect 745 -918 749 -914
rect 768 -918 772 -914
rect 823 -919 827 -915
rect 846 -919 850 -915
rect 802 -1013 806 -1009
rect 825 -1013 829 -1009
rect 1090 -1028 1094 -1024
rect 1113 -1028 1117 -1024
rect 1645 -1024 1650 -1019
rect 1660 -1024 1664 -1019
rect 1168 -1029 1172 -1025
rect 1191 -1029 1195 -1025
rect 1147 -1123 1151 -1119
rect 1170 -1123 1174 -1119
rect 755 -1162 759 -1158
rect 778 -1162 782 -1158
rect 833 -1163 837 -1159
rect 856 -1163 860 -1159
rect 812 -1257 816 -1253
rect 835 -1257 839 -1253
<< pdcontact >>
rect 672 667 676 671
rect 685 667 689 671
rect 696 667 700 671
rect 750 666 754 670
rect 763 666 767 670
rect 774 666 778 670
rect 729 572 733 576
rect 742 572 746 576
rect 753 572 757 576
rect 890 540 894 544
rect 903 540 907 544
rect 914 540 918 544
rect 968 539 972 543
rect 981 539 985 543
rect 992 539 996 543
rect 1183 502 1187 507
rect 1198 502 1202 507
rect 947 445 951 449
rect 960 445 964 449
rect 971 445 975 449
rect 685 391 689 395
rect 698 391 702 395
rect 709 391 713 395
rect 763 390 767 394
rect 776 390 780 394
rect 787 390 791 394
rect 742 296 746 300
rect 755 296 759 300
rect 766 296 770 300
rect -84 58 -80 63
rect -69 58 -65 63
rect 81 58 85 63
rect 96 58 100 63
rect 258 59 262 64
rect 273 59 277 64
rect 433 58 437 63
rect 448 58 452 63
rect 831 13 835 18
rect 846 13 850 18
rect 1079 12 1083 17
rect 1094 12 1098 17
rect 913 0 917 4
rect 922 0 926 4
rect 932 0 936 4
rect 941 0 945 4
rect 957 0 961 4
rect 966 0 970 4
rect 976 0 980 4
rect 985 0 989 4
rect 1322 21 1326 26
rect 1337 21 1341 26
rect 1161 -1 1165 3
rect 1170 -1 1174 3
rect 1180 -1 1184 3
rect 1189 -1 1193 3
rect 1205 -1 1209 3
rect 1214 -1 1218 3
rect 1224 -1 1228 3
rect 1233 -1 1237 3
rect 1591 26 1595 31
rect 1606 26 1610 31
rect 1404 8 1408 12
rect 1413 8 1417 12
rect 1423 8 1427 12
rect 1432 8 1436 12
rect 1448 8 1452 12
rect 1457 8 1461 12
rect 1467 8 1471 12
rect 1476 8 1480 12
rect 1673 13 1677 17
rect 1682 13 1686 17
rect 1692 13 1696 17
rect 1701 13 1705 17
rect 1717 13 1721 17
rect 1726 13 1730 17
rect 1736 13 1740 17
rect 1745 13 1749 17
rect 133 -55 137 -51
rect -38 -60 -34 -56
rect -25 -60 -21 -56
rect -14 -60 -10 -56
rect 19 -61 23 -56
rect 34 -61 38 -56
rect 146 -55 150 -51
rect 157 -55 161 -51
rect 190 -56 194 -51
rect 205 -56 209 -51
rect 507 -55 511 -51
rect 326 -59 330 -55
rect 339 -59 343 -55
rect 350 -59 354 -55
rect 383 -60 387 -55
rect 398 -60 402 -55
rect 520 -55 524 -51
rect 531 -55 535 -51
rect 564 -56 568 -51
rect 579 -56 583 -51
rect 1165 -116 1169 -112
rect 1178 -116 1182 -112
rect 1189 -116 1193 -112
rect 1222 -117 1226 -112
rect 1237 -117 1241 -112
rect 1541 -128 1545 -124
rect 1554 -128 1558 -124
rect 1565 -128 1569 -124
rect 1598 -129 1602 -124
rect 1613 -129 1617 -124
rect 1385 -136 1389 -132
rect 1398 -136 1402 -132
rect 1409 -136 1413 -132
rect 1442 -137 1446 -132
rect 1457 -137 1461 -132
rect 94 -199 98 -195
rect 107 -199 111 -195
rect 118 -199 122 -195
rect 151 -200 155 -195
rect 166 -200 170 -195
rect 944 -231 948 -227
rect 957 -231 961 -227
rect 968 -231 972 -227
rect 1001 -232 1005 -227
rect 1016 -232 1020 -227
rect 2095 -353 2099 -349
rect 2108 -353 2112 -349
rect 2119 -353 2123 -349
rect 2152 -354 2156 -349
rect 2167 -354 2171 -349
rect 2312 -353 2316 -349
rect 2325 -353 2329 -349
rect 2336 -353 2340 -349
rect 2369 -354 2373 -349
rect 2384 -354 2388 -349
rect 98 -397 102 -393
rect 111 -397 115 -393
rect 122 -397 126 -393
rect 155 -398 159 -393
rect 170 -398 174 -393
rect 1285 -400 1289 -396
rect 1298 -400 1302 -396
rect 1309 -400 1313 -396
rect 1342 -401 1346 -396
rect 1357 -401 1361 -396
rect 957 -417 961 -413
rect 970 -417 974 -413
rect 981 -417 985 -413
rect 1014 -418 1018 -413
rect 1029 -418 1033 -413
rect -59 -573 -55 -568
rect -44 -573 -40 -568
rect 106 -573 110 -568
rect 121 -573 125 -568
rect 283 -572 287 -567
rect 298 -572 302 -567
rect 458 -573 462 -568
rect 473 -573 477 -568
rect 158 -686 162 -682
rect -13 -691 -9 -687
rect 0 -691 4 -687
rect 11 -691 15 -687
rect 44 -692 48 -687
rect 59 -692 63 -687
rect 171 -686 175 -682
rect 182 -686 186 -682
rect 215 -687 219 -682
rect 230 -687 234 -682
rect 532 -686 536 -682
rect 351 -690 355 -686
rect 364 -690 368 -686
rect 375 -690 379 -686
rect 408 -691 412 -686
rect 423 -691 427 -686
rect 545 -686 549 -682
rect 556 -686 560 -682
rect 589 -687 593 -682
rect 604 -687 608 -682
rect 744 -887 748 -883
rect 757 -887 761 -883
rect 768 -887 772 -883
rect 822 -888 826 -884
rect 835 -888 839 -884
rect 846 -888 850 -884
rect 801 -982 805 -978
rect 814 -982 818 -978
rect 825 -982 829 -978
rect 1645 -985 1649 -980
rect 1660 -985 1664 -980
rect 1089 -997 1093 -993
rect 1102 -997 1106 -993
rect 1113 -997 1117 -993
rect 1167 -998 1171 -994
rect 1180 -998 1184 -994
rect 1191 -998 1195 -994
rect 1146 -1092 1150 -1088
rect 1159 -1092 1163 -1088
rect 1170 -1092 1174 -1088
rect 754 -1131 758 -1127
rect 767 -1131 771 -1127
rect 778 -1131 782 -1127
rect 832 -1132 836 -1128
rect 845 -1132 849 -1128
rect 856 -1132 860 -1128
rect 811 -1226 815 -1222
rect 824 -1226 828 -1222
rect 835 -1226 839 -1222
<< m2contact >>
rect 662 656 668 660
rect 741 654 748 659
rect 759 555 763 559
rect 675 380 681 384
rect 754 378 761 383
rect 959 527 966 532
rect 210 -74 214 -70
rect 833 -6 837 -2
rect 584 -74 588 -70
rect 411 -79 416 -75
rect 925 21 929 25
rect 1081 -7 1085 -3
rect 1097 -7 1102 -3
rect 1173 20 1177 24
rect 1324 2 1328 6
rect 1416 29 1420 33
rect 1593 7 1597 11
rect 1685 34 1689 38
rect 1157 -128 1161 -124
rect 172 -218 176 -214
rect 936 -243 940 -239
rect 176 -416 180 -412
rect 1021 -250 1025 -246
rect 1377 -148 1381 -144
rect 1463 -155 1467 -151
rect 610 -705 614 -701
rect 1035 -436 1039 -432
rect 1364 -420 1372 -414
rect 734 -898 740 -894
rect 813 -900 820 -895
rect 831 -999 835 -995
rect 744 -1142 750 -1138
rect 823 -1144 830 -1139
rect 1158 -1010 1165 -1005
<< nsubstratencontact >>
rect 1186 513 1190 517
rect -81 69 -77 73
rect 84 69 88 73
rect 261 70 265 74
rect 436 69 440 73
rect 834 24 838 28
rect 193 -45 197 -41
rect 567 -45 571 -41
rect 1082 23 1086 27
rect 1325 32 1329 36
rect 1594 37 1598 41
rect 22 -50 26 -46
rect 386 -49 390 -45
rect 1225 -106 1229 -102
rect 1601 -118 1605 -114
rect 1445 -126 1449 -122
rect 154 -189 158 -185
rect 1004 -221 1008 -217
rect 2155 -343 2159 -339
rect 2372 -343 2376 -339
rect 158 -387 162 -383
rect 1345 -390 1349 -386
rect 1017 -407 1021 -403
rect -56 -562 -52 -558
rect 109 -562 113 -558
rect 286 -561 290 -557
rect 461 -562 465 -558
rect 218 -676 222 -672
rect 592 -676 596 -672
rect 47 -681 51 -677
rect 411 -680 415 -676
rect 1648 -974 1652 -970
<< labels >>
rlabel metal1 -71 71 -71 71 5 vdd
rlabel metal1 -76 9 -76 9 1 gnd
rlabel metal1 -78 41 -78 41 1 A0
rlabel metal1 -67 41 -67 41 1 na0
rlabel metal1 94 71 94 71 5 vdd
rlabel metal1 89 9 89 9 1 gnd
rlabel metal1 87 41 87 41 1 A1
rlabel metal1 98 41 98 41 1 na1
rlabel metal1 -1 -49 -1 -49 1 vdd
rlabel metal1 2 -104 2 -104 1 gnd
rlabel metal1 -37 -77 -37 -77 1 B0
rlabel metal1 38 -77 38 -77 1 w7
rlabel metal1 170 -44 170 -44 1 vdd
rlabel metal1 173 -99 173 -99 1 gnd
rlabel metal1 134 -72 134 -72 1 B1
rlabel metal1 208 -73 208 -73 1 w5
rlabel metal1 446 71 446 71 5 vdd
rlabel metal1 441 9 441 9 1 gnd
rlabel metal1 439 41 439 41 1 A3
rlabel metal1 450 40 450 40 1 na3
rlabel metal1 544 -44 544 -44 1 vdd
rlabel metal1 547 -99 547 -99 1 gnd
rlabel metal1 510 -72 510 -72 1 B3
rlabel metal1 584 -73 584 -73 1 w1
rlabel metal1 401 -76 401 -76 1 w3
rlabel metal1 328 -75 328 -75 1 B2
rlabel metal1 366 -103 366 -103 1 gnd
rlabel metal1 363 -48 363 -48 1 vdd
rlabel metal1 275 41 275 41 1 na2
rlabel metal1 263 42 263 42 1 A2
rlabel metal1 266 10 266 10 1 gnd
rlabel metal1 271 72 271 72 5 vdd
rlabel metal1 970 -36 970 -36 1 gnd
rlabel metal1 969 17 969 17 1 vdd
rlabel metal1 844 26 844 26 5 vdd
rlabel metal1 839 -36 839 -36 1 gnd
rlabel metal1 953 -14 953 -14 1 A3
rlabel polysilicon 982 -15 982 -15 1 B3
rlabel metal1 849 -6 849 -6 1 x3
rlabel metal1 1218 -37 1218 -37 1 gnd
rlabel metal1 1217 16 1217 16 1 vdd
rlabel metal1 1092 25 1092 25 5 vdd
rlabel metal1 1087 -37 1087 -37 1 gnd
rlabel metal1 1200 -14 1200 -14 1 A2
rlabel polysilicon 1230 -15 1230 -15 1 B2
rlabel metal1 1096 -6 1096 -6 1 x2
rlabel metal1 1461 -28 1461 -28 1 gnd
rlabel metal1 1460 25 1460 25 1 vdd
rlabel metal1 1335 34 1335 34 5 vdd
rlabel metal1 1330 -28 1330 -28 1 gnd
rlabel metal1 1442 -5 1442 -5 1 A1
rlabel polysilicon 1473 -7 1473 -7 1 B1
rlabel metal1 1339 2 1339 2 1 x1
rlabel metal1 1599 -23 1599 -23 1 gnd
rlabel metal1 1604 39 1604 39 5 vdd
rlabel metal1 1729 30 1729 30 1 vdd
rlabel metal1 1730 -23 1730 -23 1 gnd
rlabel metal1 1609 7 1609 7 1 x0
rlabel metal1 1710 1 1710 1 1 A0
rlabel polysilicon 1742 -2 1742 -2 1 B0
rlabel metal1 -46 -560 -46 -560 5 vdd
rlabel metal1 -51 -622 -51 -622 1 gnd
rlabel metal1 119 -560 119 -560 5 vdd
rlabel metal1 114 -622 114 -622 1 gnd
rlabel metal1 24 -680 24 -680 1 vdd
rlabel metal1 27 -735 27 -735 1 gnd
rlabel metal1 195 -675 195 -675 1 vdd
rlabel metal1 198 -730 198 -730 1 gnd
rlabel metal1 471 -560 471 -560 5 vdd
rlabel metal1 466 -622 466 -622 1 gnd
rlabel metal1 569 -675 569 -675 1 vdd
rlabel metal1 572 -730 572 -730 1 gnd
rlabel metal1 391 -734 391 -734 1 gnd
rlabel metal1 388 -679 388 -679 1 vdd
rlabel metal1 291 -621 291 -621 1 gnd
rlabel metal1 296 -559 296 -559 5 vdd
rlabel metal1 -53 -589 -53 -589 1 B0
rlabel metal1 -41 -589 -41 -589 1 nb0
rlabel metal1 112 -589 112 -589 1 B1
rlabel metal1 129 -589 129 -589 1 nb1
rlabel metal1 288 -589 288 -589 1 B2
rlabel metal1 304 -588 304 -588 1 nb2
rlabel metal1 463 -590 463 -590 1 B3
rlabel metal1 479 -590 479 -590 1 nb3
rlabel metal1 -14 -708 -14 -708 1 A0
rlabel metal1 64 -708 64 -708 1 w8
rlabel metal1 159 -703 159 -703 1 A1
rlabel metal1 350 -707 350 -707 1 A2
rlabel metal1 428 -707 428 -707 1 w4
rlabel metal1 533 -703 533 -703 1 A3
rlabel metal1 608 -703 608 -703 1 w2
rlabel metal1 983 -218 983 -218 1 vdd
rlabel metal1 983 -272 983 -272 1 gnd
rlabel metal1 1020 -248 1020 -248 1 t1
rlabel metal1 996 -404 996 -404 1 vdd
rlabel metal1 996 -458 996 -458 1 gnd
rlabel metal1 1034 -434 1034 -434 1 t2
rlabel metal1 1204 -103 1204 -103 1 vdd
rlabel metal1 1204 -157 1204 -157 1 gnd
rlabel metal1 1240 -133 1240 -133 1 o1
rlabel metal1 1424 -177 1424 -177 1 gnd
rlabel metal1 1424 -123 1424 -123 1 vdd
rlabel metal1 1461 -153 1461 -153 1 t3
rlabel metal1 1324 -441 1324 -441 1 gnd
rlabel metal1 1324 -387 1324 -387 1 vdd
rlabel metal1 235 -703 235 -703 1 w6
rlabel metal1 1361 -418 1361 -418 1 t4
rlabel metal1 1580 -169 1580 -169 1 gnd
rlabel metal1 1580 -115 1580 -115 1 vdd
rlabel metal1 1618 -146 1618 -146 1 o2
rlabel metal1 133 -240 133 -240 1 gnd
rlabel metal1 133 -186 133 -186 1 vdd
rlabel metal1 137 -438 137 -438 1 gnd
rlabel metal1 137 -384 137 -384 1 vdd
rlabel metal1 170 -217 170 -217 1 t5
rlabel metal1 176 -414 176 -414 1 t6
rlabel metal1 737 402 737 402 5 vdd
rlabel metal1 755 309 755 309 1 vdd
rlabel metal1 698 348 698 348 1 gnd
rlabel metal1 778 347 778 347 1 gnd
rlabel metal1 757 253 757 253 1 gnd
rlabel metal1 772 280 772 280 1 l1
rlabel metal1 724 678 724 678 5 vdd
rlabel metal1 742 585 742 585 1 vdd
rlabel metal1 685 624 685 624 1 gnd
rlabel metal1 765 623 765 623 1 gnd
rlabel metal1 744 529 744 529 1 gnd
rlabel metal1 758 557 758 557 1 l2
rlabel metal1 942 551 942 551 5 vdd
rlabel metal1 960 458 960 458 1 vdd
rlabel metal1 903 497 903 497 1 gnd
rlabel metal1 962 402 962 402 1 gnd
rlabel metal1 978 431 978 431 1 y0
rlabel metal1 983 496 983 496 1 gnd
rlabel metal1 796 -876 796 -876 5 vdd
rlabel metal1 814 -969 814 -969 1 vdd
rlabel metal1 757 -930 757 -930 1 gnd
rlabel metal1 837 -931 837 -931 1 gnd
rlabel metal1 816 -1025 816 -1025 1 gnd
rlabel metal1 829 -997 829 -997 1 g1
rlabel metal1 806 -1120 806 -1120 5 vdd
rlabel metal1 824 -1213 824 -1213 1 vdd
rlabel metal1 767 -1174 767 -1174 1 gnd
rlabel metal1 847 -1175 847 -1175 1 gnd
rlabel metal1 826 -1269 826 -1269 1 gnd
rlabel metal1 1141 -986 1141 -986 5 vdd
rlabel metal1 1159 -1079 1159 -1079 1 vdd
rlabel metal1 1102 -1040 1102 -1040 1 gnd
rlabel metal1 1182 -1041 1182 -1041 1 gnd
rlabel metal1 1161 -1135 1161 -1135 1 gnd
rlabel metal1 1174 -1108 1174 -1107 1 y1
rlabel metal1 838 -1241 838 -1241 1 g2
rlabel metal1 1191 453 1191 453 1 gnd
rlabel metal1 1196 515 1196 515 5 vdd
rlabel metal1 1200 484 1200 484 1 y0d
rlabel metal1 1653 -1034 1653 -1034 1 gnd
rlabel metal1 1658 -972 1658 -972 5 vdd
rlabel metal1 1663 -1003 1663 -1003 1 y1d
rlabel metal1 2134 -394 2134 -394 1 gnd
rlabel metal1 2134 -340 2134 -340 1 vdd
rlabel metal1 2171 -371 2171 -371 1 e1
rlabel metal1 2351 -394 2351 -394 1 gnd
rlabel metal1 2351 -340 2351 -340 1 vdd
rlabel metal1 2388 -371 2388 -371 1 y2
rlabel metal1 2310 -363 2310 -363 1 D2
<< end >>
