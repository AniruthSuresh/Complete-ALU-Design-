magic
tech scmos
timestamp 1699698287
<< checkpaint >>
rect -66 -4 0 82
<< metal1 >>
rect -20 63 1 67
rect 41 63 42 67
rect -50 42 -44 46
rect -50 34 -45 38
rect -20 37 -19 38
rect -20 33 16 37
rect 28 35 31 37
rect 29 34 31 35
rect -18 9 0 13
rect -18 8 10 9
rect -18 5 12 8
use nand2  nand2_0
timestamp 1699617909
transform 1 0 -45 0 1 33
box -7 -23 31 35
use not  not_0
timestamp 1699617317
transform 1 0 21 0 1 34
box -21 -34 21 33
<< labels >>
rlabel metal1 -50 44 -50 44 3 A
rlabel metal1 -50 36 -50 36 3 B
rlabel metal1 42 65 42 65 6 vdd
rlabel metal1 6 9 6 9 1 gnd
rlabel metal1 31 36 31 36 1 out
<< end >>
