
.subckt AND node_a node_b node_out vdd gnd

	X1 node_a node_b node_c vdd gnd NAND
	X2 node_c node_c node_out vdd gnd NAND

.ends AND

